module pla_lined (
	movEa,
	col,
	opcode,
	lineBmap,
	palIll,
	plaA1,
	plaA2,
	plaA3
);
	reg _sv2v_0;
	input [3:0] movEa;
	input [3:0] col;
	input [15:0] opcode;
	input [15:0] lineBmap;
	output wire palIll;
	output wire [9:0] plaA1;
	output wire [9:0] plaA2;
	output wire [9:0] plaA3;
	wire [3:0] line = opcode[15:12];
	wire [2:0] row86 = opcode[8:6];
	reg [15:0] arIll;
	reg [9:0] arA1 [15:0];
	reg [9:0] arA23 [15:0];
	reg [9:0] scA3;
	reg illMisc;
	reg [9:0] a1Misc;
	assign palIll = |(arIll & lineBmap);
	assign plaA1 = arA1[line];
	assign plaA2 = arA23[line];
	assign plaA3 = (lineBmap[0] ? scA3 : arA23[line]);
	always @(*) begin
		if (_sv2v_0)
			;
		arIll['h6] = 1'b0;
		arA23['h6] = 1'sbx;
		if (opcode[11:8] == 4'h1)
			arA1['h6] = (|opcode[7:0] ? 'h89 : 'ha9);
		else
			arA1['h6] = (|opcode[7:0] ? 'h308 : 'h68);
		arIll['h7] = opcode[8];
		arA23['h7] = 1'sbx;
		arA1['h7] = 'h23b;
		arIll['ha] = 1'b1;
		arIll['hf] = 1'b1;
		arA1['ha] = 1'sbx;
		arA1['hf] = 1'sbx;
		arA23['ha] = 1'sbx;
		arA23['hf] = 1'sbx;
	end
	always @(*) begin
		if (_sv2v_0)
			;
		if ((~opcode[11] & opcode[7]) & opcode[6]) begin
			arA23['he] = 'h3c7;
			(* full_case, parallel_case *)
			case (col)
				2: begin
					arIll['he] = 1'b0;
					arA1['he] = 'h6;
				end
				3: begin
					arIll['he] = 1'b0;
					arA1['he] = 'h21c;
				end
				4: begin
					arIll['he] = 1'b0;
					arA1['he] = 'h103;
				end
				5: begin
					arIll['he] = 1'b0;
					arA1['he] = 'h1c2;
				end
				6: begin
					arIll['he] = 1'b0;
					arA1['he] = 'h1e3;
				end
				7: begin
					arIll['he] = 1'b0;
					arA1['he] = 'ha;
				end
				8: begin
					arIll['he] = 1'b0;
					arA1['he] = 'h1e2;
				end
				default: begin
					arIll['he] = 1'b1;
					arA1['he] = 1'sbx;
				end
			endcase
		end
		else begin
			arA23['he] = 1'sbx;
			(* full_case, parallel_case *)
			case (opcode[7:6])
				2'b00, 2'b01: begin
					arIll['he] = 1'b0;
					arA1['he] = (opcode[5] ? 'h382 : 'h381);
				end
				2'b10: begin
					arIll['he] = 1'b0;
					arA1['he] = (opcode[5] ? 'h386 : 'h385);
				end
				2'b11: begin
					arIll['he] = 1'b1;
					arA1['he] = 1'sbx;
				end
			endcase
		end
	end
	always @(*) begin
		if (_sv2v_0)
			;
		illMisc = 1'b0;
		case (opcode[5:3])
			3'b000, 3'b001: a1Misc = 'h1d0;
			3'b010: a1Misc = 'h30b;
			3'b011: a1Misc = 'h119;
			3'b100: a1Misc = 'h2f5;
			3'b101: a1Misc = 'h230;
			3'b110:
				case (opcode[2:0])
					3'b110: a1Misc = 'h6d;
					3'b000: a1Misc = 'h3a6;
					3'b001: a1Misc = 'h363;
					3'b010: a1Misc = 'h3a2;
					3'b011: a1Misc = 'h12a;
					3'b111: a1Misc = 'h12a;
					3'b101: a1Misc = 'h126;
					default: begin
						illMisc = 1'b1;
						a1Misc = 1'sbx;
					end
				endcase
			default: begin
				illMisc = 1'b1;
				a1Misc = 1'sbx;
			end
		endcase
	end
	always @(*) begin
		if (_sv2v_0)
			;
		if ((opcode[11:6] & 'h1f) == 'h8)
			(* full_case, parallel_case *)
			case (col)
				0: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h100;
					scA3 = 1'sbx;
				end
				1: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				2: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h6;
					scA3 = 'h299;
				end
				3: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h21c;
					scA3 = 'h299;
				end
				4: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h103;
					scA3 = 'h299;
				end
				5: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h1c2;
					scA3 = 'h299;
				end
				6: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h1e3;
					scA3 = 'h299;
				end
				7: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'ha;
					scA3 = 'h299;
				end
				8: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h1e2;
					scA3 = 'h299;
				end
				9: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				10: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				11: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h1cc;
					scA3 = 1'sbx;
				end
				default: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
			endcase
		else if ((opcode[11:6] & 'h37) == 'h0)
			(* full_case, parallel_case *)
			case (col)
				0: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h100;
					scA3 = 1'sbx;
				end
				1: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				2: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h6;
					scA3 = 'h299;
				end
				3: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h21c;
					scA3 = 'h299;
				end
				4: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h103;
					scA3 = 'h299;
				end
				5: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h1c2;
					scA3 = 'h299;
				end
				6: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h1e3;
					scA3 = 'h299;
				end
				7: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'ha;
					scA3 = 'h299;
				end
				8: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h1e2;
					scA3 = 'h299;
				end
				9: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				10: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				11: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h1cc;
					scA3 = 1'sbx;
				end
				default: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
			endcase
		else if ((opcode[11:6] & 'h1f) == 'h9)
			(* full_case, parallel_case *)
			case (col)
				0: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h100;
					scA3 = 1'sbx;
				end
				1: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				2: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h6;
					scA3 = 'h299;
				end
				3: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h21c;
					scA3 = 'h299;
				end
				4: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h103;
					scA3 = 'h299;
				end
				5: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h1c2;
					scA3 = 'h299;
				end
				6: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h1e3;
					scA3 = 'h299;
				end
				7: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'ha;
					scA3 = 'h299;
				end
				8: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h1e2;
					scA3 = 'h299;
				end
				9: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				10: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				11: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h1cc;
					scA3 = 1'sbx;
				end
				default: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
			endcase
		else if ((opcode[11:6] & 'h37) == 'h1)
			(* full_case, parallel_case *)
			case (col)
				0: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h100;
					scA3 = 1'sbx;
				end
				1: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				2: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h6;
					scA3 = 'h299;
				end
				3: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h21c;
					scA3 = 'h299;
				end
				4: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h103;
					scA3 = 'h299;
				end
				5: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h1c2;
					scA3 = 'h299;
				end
				6: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h1e3;
					scA3 = 'h299;
				end
				7: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'ha;
					scA3 = 'h299;
				end
				8: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h1e2;
					scA3 = 'h299;
				end
				9: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				10: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				11: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h1cc;
					scA3 = 1'sbx;
				end
				default: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
			endcase
		else if ((opcode[11:6] & 'h1f) == 'ha)
			(* full_case, parallel_case *)
			case (col)
				0: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h3e0;
					arA23['h0] = 'h10c;
					scA3 = 1'sbx;
				end
				1: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				2: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h3e0;
					arA23['h0] = 'hb;
					scA3 = 'h29d;
				end
				3: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h3e0;
					arA23['h0] = 'hf;
					scA3 = 'h29d;
				end
				4: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h3e0;
					arA23['h0] = 'h179;
					scA3 = 'h29d;
				end
				5: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h3e0;
					arA23['h0] = 'h1c6;
					scA3 = 'h29d;
				end
				6: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h3e0;
					arA23['h0] = 'h1e7;
					scA3 = 'h29d;
				end
				7: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h3e0;
					arA23['h0] = 'he;
					scA3 = 'h29d;
				end
				8: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h3e0;
					arA23['h0] = 'h1e6;
					scA3 = 'h29d;
				end
				9: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				10: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				11: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				default: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
			endcase
		else if ((opcode[11:6] & 'h37) == 'h2)
			(* full_case, parallel_case *)
			case (col)
				0: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h3e0;
					arA23['h0] = 'h10c;
					scA3 = 1'sbx;
				end
				1: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				2: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h3e0;
					arA23['h0] = 'hb;
					scA3 = 'h29d;
				end
				3: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h3e0;
					arA23['h0] = 'hf;
					scA3 = 'h29d;
				end
				4: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h3e0;
					arA23['h0] = 'h179;
					scA3 = 'h29d;
				end
				5: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h3e0;
					arA23['h0] = 'h1c6;
					scA3 = 'h29d;
				end
				6: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h3e0;
					arA23['h0] = 'h1e7;
					scA3 = 'h29d;
				end
				7: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h3e0;
					arA23['h0] = 'he;
					scA3 = 'h29d;
				end
				8: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h3e0;
					arA23['h0] = 'h1e6;
					scA3 = 'h29d;
				end
				9: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				10: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				11: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				default: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
			endcase
		else if ((opcode[11:6] & 'h37) == 'h10)
			(* full_case, parallel_case *)
			case (col)
				0: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h100;
					scA3 = 1'sbx;
				end
				1: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				2: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h6;
					scA3 = 'h299;
				end
				3: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h21c;
					scA3 = 'h299;
				end
				4: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h103;
					scA3 = 'h299;
				end
				5: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h1c2;
					scA3 = 'h299;
				end
				6: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h1e3;
					scA3 = 'h299;
				end
				7: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'ha;
					scA3 = 'h299;
				end
				8: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h1e2;
					scA3 = 'h299;
				end
				9: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				10: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				11: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				default: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
			endcase
		else if ((opcode[11:6] & 'h37) == 'h11)
			(* full_case, parallel_case *)
			case (col)
				0: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h100;
					scA3 = 1'sbx;
				end
				1: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				2: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h6;
					scA3 = 'h299;
				end
				3: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h21c;
					scA3 = 'h299;
				end
				4: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h103;
					scA3 = 'h299;
				end
				5: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h1c2;
					scA3 = 'h299;
				end
				6: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h1e3;
					scA3 = 'h299;
				end
				7: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'ha;
					scA3 = 'h299;
				end
				8: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h1e2;
					scA3 = 'h299;
				end
				9: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				10: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				11: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				default: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
			endcase
		else if ((opcode[11:6] & 'h37) == 'h12)
			(* full_case, parallel_case *)
			case (col)
				0: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h3e0;
					arA23['h0] = 'h10c;
					scA3 = 1'sbx;
				end
				1: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				2: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h3e0;
					arA23['h0] = 'hb;
					scA3 = 'h29d;
				end
				3: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h3e0;
					arA23['h0] = 'hf;
					scA3 = 'h29d;
				end
				4: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h3e0;
					arA23['h0] = 'h179;
					scA3 = 'h29d;
				end
				5: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h3e0;
					arA23['h0] = 'h1c6;
					scA3 = 'h29d;
				end
				6: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h3e0;
					arA23['h0] = 'h1e7;
					scA3 = 'h29d;
				end
				7: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h3e0;
					arA23['h0] = 'he;
					scA3 = 'h29d;
				end
				8: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h3e0;
					arA23['h0] = 'h1e6;
					scA3 = 'h29d;
				end
				9: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				10: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				11: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				default: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
			endcase
		else if ((opcode[11:6] & 'h7) == 'h4)
			(* full_case, parallel_case *)
			case (col)
				0: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h3e7;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				1: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h1d2;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				2: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h6;
					arA23['h0] = 1'sbx;
					scA3 = 'h215;
				end
				3: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h21c;
					arA23['h0] = 1'sbx;
					scA3 = 'h215;
				end
				4: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h103;
					arA23['h0] = 1'sbx;
					scA3 = 'h215;
				end
				5: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h1c2;
					arA23['h0] = 1'sbx;
					scA3 = 'h215;
				end
				6: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h1e3;
					arA23['h0] = 1'sbx;
					scA3 = 'h215;
				end
				7: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'ha;
					arA23['h0] = 1'sbx;
					scA3 = 'h215;
				end
				8: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h1e2;
					arA23['h0] = 1'sbx;
					scA3 = 'h215;
				end
				9: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h1c2;
					arA23['h0] = 1'sbx;
					scA3 = 'h215;
				end
				10: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h1e3;
					arA23['h0] = 1'sbx;
					scA3 = 'h215;
				end
				11: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'hea;
					arA23['h0] = 'hab;
					scA3 = 1'sbx;
				end
				default: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
			endcase
		else if ((opcode[11:6] & 'h7) == 'h5)
			(* full_case, parallel_case *)
			case (col)
				0: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h3ef;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				1: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h1d6;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				2: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h6;
					arA23['h0] = 1'sbx;
					scA3 = 'h81;
				end
				3: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h21c;
					arA23['h0] = 1'sbx;
					scA3 = 'h81;
				end
				4: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h103;
					arA23['h0] = 1'sbx;
					scA3 = 'h81;
				end
				5: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h1c2;
					arA23['h0] = 1'sbx;
					scA3 = 'h81;
				end
				6: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h1e3;
					arA23['h0] = 1'sbx;
					scA3 = 'h81;
				end
				7: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'ha;
					arA23['h0] = 1'sbx;
					scA3 = 'h81;
				end
				8: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h1e2;
					arA23['h0] = 1'sbx;
					scA3 = 'h81;
				end
				9: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				10: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				11: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				default: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
			endcase
		else if ((opcode[11:6] & 'h7) == 'h7)
			(* full_case, parallel_case *)
			case (col)
				0: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h3ef;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				1: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h1ce;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				2: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h6;
					arA23['h0] = 1'sbx;
					scA3 = 'h81;
				end
				3: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h21c;
					arA23['h0] = 1'sbx;
					scA3 = 'h81;
				end
				4: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h103;
					arA23['h0] = 1'sbx;
					scA3 = 'h81;
				end
				5: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h1c2;
					arA23['h0] = 1'sbx;
					scA3 = 'h81;
				end
				6: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h1e3;
					arA23['h0] = 1'sbx;
					scA3 = 'h81;
				end
				7: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'ha;
					arA23['h0] = 1'sbx;
					scA3 = 'h81;
				end
				8: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h1e2;
					arA23['h0] = 1'sbx;
					scA3 = 'h81;
				end
				9: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				10: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				11: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				default: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
			endcase
		else if ((opcode[11:6] & 'h7) == 'h6)
			(* full_case, parallel_case *)
			case (col)
				0: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h3eb;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				1: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h1ca;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				2: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h6;
					arA23['h0] = 1'sbx;
					scA3 = 'h69;
				end
				3: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h21c;
					arA23['h0] = 1'sbx;
					scA3 = 'h69;
				end
				4: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h103;
					arA23['h0] = 1'sbx;
					scA3 = 'h69;
				end
				5: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h1c2;
					arA23['h0] = 1'sbx;
					scA3 = 'h69;
				end
				6: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h1e3;
					arA23['h0] = 1'sbx;
					scA3 = 'h69;
				end
				7: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'ha;
					arA23['h0] = 1'sbx;
					scA3 = 'h69;
				end
				8: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h1e2;
					arA23['h0] = 1'sbx;
					scA3 = 'h69;
				end
				9: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				10: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				11: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				default: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
			endcase
		else if (opcode[11:6] == 'h20)
			(* full_case, parallel_case *)
			case (col)
				0: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h3e7;
					scA3 = 1'sbx;
				end
				1: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				2: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h6;
					scA3 = 'h215;
				end
				3: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h21c;
					scA3 = 'h215;
				end
				4: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h103;
					scA3 = 'h215;
				end
				5: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h1c2;
					scA3 = 'h215;
				end
				6: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h1e3;
					scA3 = 'h215;
				end
				7: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'ha;
					scA3 = 'h215;
				end
				8: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h1e2;
					scA3 = 'h215;
				end
				9: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h1c2;
					scA3 = 'h215;
				end
				10: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h1e3;
					scA3 = 'h215;
				end
				11: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				default: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
			endcase
		else if (opcode[11:6] == 'h21)
			(* full_case, parallel_case *)
			case (col)
				0: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h3ef;
					scA3 = 1'sbx;
				end
				1: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				2: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h6;
					scA3 = 'h81;
				end
				3: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h21c;
					scA3 = 'h81;
				end
				4: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h103;
					scA3 = 'h81;
				end
				5: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h1c2;
					scA3 = 'h81;
				end
				6: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h1e3;
					scA3 = 'h81;
				end
				7: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'ha;
					scA3 = 'h81;
				end
				8: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h1e2;
					scA3 = 'h81;
				end
				9: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				10: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				11: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				default: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
			endcase
		else if (opcode[11:6] == 'h23)
			(* full_case, parallel_case *)
			case (col)
				0: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h3ef;
					scA3 = 1'sbx;
				end
				1: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				2: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h6;
					scA3 = 'h81;
				end
				3: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h21c;
					scA3 = 'h81;
				end
				4: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h103;
					scA3 = 'h81;
				end
				5: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h1c2;
					scA3 = 'h81;
				end
				6: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h1e3;
					scA3 = 'h81;
				end
				7: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'ha;
					scA3 = 'h81;
				end
				8: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h1e2;
					scA3 = 'h81;
				end
				9: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				10: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				11: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				default: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
			endcase
		else if (opcode[11:6] == 'h22)
			(* full_case, parallel_case *)
			case (col)
				0: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h3eb;
					scA3 = 1'sbx;
				end
				1: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				2: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h6;
					scA3 = 'h69;
				end
				3: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h21c;
					scA3 = 'h69;
				end
				4: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h103;
					scA3 = 'h69;
				end
				5: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h1c2;
					scA3 = 'h69;
				end
				6: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h1e3;
					scA3 = 'h69;
				end
				7: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'ha;
					scA3 = 'h69;
				end
				8: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h1e2;
					scA3 = 'h69;
				end
				9: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				10: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				11: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				default: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
			endcase
		else if (opcode[11:6] == 'h30)
			(* full_case, parallel_case *)
			case (col)
				0: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h108;
					scA3 = 1'sbx;
				end
				1: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				2: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h6;
					scA3 = 'h87;
				end
				3: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h21c;
					scA3 = 'h87;
				end
				4: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h103;
					scA3 = 'h87;
				end
				5: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h1c2;
					scA3 = 'h87;
				end
				6: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h1e3;
					scA3 = 'h87;
				end
				7: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'ha;
					scA3 = 'h87;
				end
				8: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h1e2;
					scA3 = 'h87;
				end
				9: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				10: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				11: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				default: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
			endcase
		else if (opcode[11:6] == 'h31)
			(* full_case, parallel_case *)
			case (col)
				0: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h108;
					scA3 = 1'sbx;
				end
				1: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				2: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h6;
					scA3 = 'h87;
				end
				3: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h21c;
					scA3 = 'h87;
				end
				4: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h103;
					scA3 = 'h87;
				end
				5: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h1c2;
					scA3 = 'h87;
				end
				6: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h1e3;
					scA3 = 'h87;
				end
				7: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'ha;
					scA3 = 'h87;
				end
				8: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h2b9;
					arA23['h0] = 'h1e2;
					scA3 = 'h87;
				end
				9: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				10: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				11: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				default: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
			endcase
		else if (opcode[11:6] == 'h32)
			(* full_case, parallel_case *)
			case (col)
				0: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h3e0;
					arA23['h0] = 'h104;
					scA3 = 1'sbx;
				end
				1: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				2: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h3e0;
					arA23['h0] = 'hb;
					scA3 = 'h8f;
				end
				3: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h3e0;
					arA23['h0] = 'hf;
					scA3 = 'h8f;
				end
				4: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h3e0;
					arA23['h0] = 'h179;
					scA3 = 'h8f;
				end
				5: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h3e0;
					arA23['h0] = 'h1c6;
					scA3 = 'h8f;
				end
				6: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h3e0;
					arA23['h0] = 'h1e7;
					scA3 = 'h8f;
				end
				7: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h3e0;
					arA23['h0] = 'he;
					scA3 = 'h8f;
				end
				8: begin
					arIll['h0] = 1'b0;
					arA1['h0] = 'h3e0;
					arA23['h0] = 'h1e6;
					scA3 = 'h8f;
				end
				9: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				10: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				11: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
				default: begin
					arIll['h0] = 1'b1;
					arA1['h0] = 1'sbx;
					arA23['h0] = 1'sbx;
					scA3 = 1'sbx;
				end
			endcase
		else begin
			arIll['h0] = 1'b1;
			arA1['h0] = 1'sbx;
			arA23['h0] = 1'sbx;
			scA3 = 1'sbx;
		end
	end
	always @(*) begin
		if (_sv2v_0)
			;
		if ((opcode[11:6] & 'h27) == 'h0)
			(* full_case, parallel_case *)
			case (col)
				0: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h133;
					arA23['h4] = 1'sbx;
				end
				1: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				2: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h6;
					arA23['h4] = 'h2b8;
				end
				3: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h21c;
					arA23['h4] = 'h2b8;
				end
				4: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h103;
					arA23['h4] = 'h2b8;
				end
				5: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1c2;
					arA23['h4] = 'h2b8;
				end
				6: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1e3;
					arA23['h4] = 'h2b8;
				end
				7: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'ha;
					arA23['h4] = 'h2b8;
				end
				8: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1e2;
					arA23['h4] = 'h2b8;
				end
				9: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				10: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				11: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				default: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
			endcase
		else if ((opcode[11:6] & 'h27) == 'h1)
			(* full_case, parallel_case *)
			case (col)
				0: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h133;
					arA23['h4] = 1'sbx;
				end
				1: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				2: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h6;
					arA23['h4] = 'h2b8;
				end
				3: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h21c;
					arA23['h4] = 'h2b8;
				end
				4: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h103;
					arA23['h4] = 'h2b8;
				end
				5: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1c2;
					arA23['h4] = 'h2b8;
				end
				6: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1e3;
					arA23['h4] = 'h2b8;
				end
				7: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'ha;
					arA23['h4] = 'h2b8;
				end
				8: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1e2;
					arA23['h4] = 'h2b8;
				end
				9: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				10: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				11: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				default: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
			endcase
		else if ((opcode[11:6] & 'h27) == 'h2)
			(* full_case, parallel_case *)
			case (col)
				0: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h137;
					arA23['h4] = 1'sbx;
				end
				1: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				2: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'hb;
					arA23['h4] = 'h2bc;
				end
				3: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'hf;
					arA23['h4] = 'h2bc;
				end
				4: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h179;
					arA23['h4] = 'h2bc;
				end
				5: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1c6;
					arA23['h4] = 'h2bc;
				end
				6: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1e7;
					arA23['h4] = 'h2bc;
				end
				7: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'he;
					arA23['h4] = 'h2bc;
				end
				8: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1e6;
					arA23['h4] = 'h2bc;
				end
				9: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				10: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				11: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				default: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
			endcase
		else if (opcode[11:6] == 'h3)
			(* full_case, parallel_case *)
			case (col)
				0: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h3a5;
					arA23['h4] = 1'sbx;
				end
				1: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				2: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h6;
					arA23['h4] = 'h3a1;
				end
				3: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h21c;
					arA23['h4] = 'h3a1;
				end
				4: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h103;
					arA23['h4] = 'h3a1;
				end
				5: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1c2;
					arA23['h4] = 'h3a1;
				end
				6: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1e3;
					arA23['h4] = 'h3a1;
				end
				7: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'ha;
					arA23['h4] = 'h3a1;
				end
				8: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1e2;
					arA23['h4] = 'h3a1;
				end
				9: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				10: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				11: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				default: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
			endcase
		else if (opcode[11:6] == 'h13)
			(* full_case, parallel_case *)
			case (col)
				0: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h301;
					arA23['h4] = 1'sbx;
				end
				1: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				2: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h6;
					arA23['h4] = 'h159;
				end
				3: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h21c;
					arA23['h4] = 'h159;
				end
				4: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h103;
					arA23['h4] = 'h159;
				end
				5: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1c2;
					arA23['h4] = 'h159;
				end
				6: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1e3;
					arA23['h4] = 'h159;
				end
				7: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'ha;
					arA23['h4] = 'h159;
				end
				8: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1e2;
					arA23['h4] = 'h159;
				end
				9: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1c2;
					arA23['h4] = 'h159;
				end
				10: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1e3;
					arA23['h4] = 'h159;
				end
				11: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'hea;
					arA23['h4] = 'h301;
				end
				default: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
			endcase
		else if (opcode[11:6] == 'h1b)
			(* full_case, parallel_case *)
			case (col)
				0: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h301;
					arA23['h4] = 1'sbx;
				end
				1: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				2: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h6;
					arA23['h4] = 'h159;
				end
				3: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h21c;
					arA23['h4] = 'h159;
				end
				4: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h103;
					arA23['h4] = 'h159;
				end
				5: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1c2;
					arA23['h4] = 'h159;
				end
				6: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1e3;
					arA23['h4] = 'h159;
				end
				7: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'ha;
					arA23['h4] = 'h159;
				end
				8: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1e2;
					arA23['h4] = 'h159;
				end
				9: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1c2;
					arA23['h4] = 'h159;
				end
				10: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1e3;
					arA23['h4] = 'h159;
				end
				11: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'hea;
					arA23['h4] = 'h301;
				end
				default: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
			endcase
		else if (opcode[11:6] == 'h20)
			(* full_case, parallel_case *)
			case (col)
				0: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h13b;
					arA23['h4] = 1'sbx;
				end
				1: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				2: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h6;
					arA23['h4] = 'h15c;
				end
				3: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h21c;
					arA23['h4] = 'h15c;
				end
				4: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h103;
					arA23['h4] = 'h15c;
				end
				5: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1c2;
					arA23['h4] = 'h15c;
				end
				6: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1e3;
					arA23['h4] = 'h15c;
				end
				7: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'ha;
					arA23['h4] = 'h15c;
				end
				8: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1e2;
					arA23['h4] = 'h15c;
				end
				9: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				10: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				11: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				default: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
			endcase
		else if (opcode[11:6] == 'h21)
			(* full_case, parallel_case *)
			case (col)
				0: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h341;
					arA23['h4] = 1'sbx;
				end
				1: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				2: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h17c;
					arA23['h4] = 1'sbx;
				end
				3: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				4: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				5: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h17d;
					arA23['h4] = 1'sbx;
				end
				6: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1ff;
					arA23['h4] = 1'sbx;
				end
				7: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h178;
					arA23['h4] = 1'sbx;
				end
				8: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1fa;
					arA23['h4] = 1'sbx;
				end
				9: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h17d;
					arA23['h4] = 1'sbx;
				end
				10: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1ff;
					arA23['h4] = 1'sbx;
				end
				11: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				default: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
			endcase
		else if (opcode[11:6] == 'h22)
			(* full_case, parallel_case *)
			case (col)
				0: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h133;
					arA23['h4] = 1'sbx;
				end
				1: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				2: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h3a0;
					arA23['h4] = 1'sbx;
				end
				3: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				4: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h3a4;
					arA23['h4] = 1'sbx;
				end
				5: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1f1;
					arA23['h4] = 1'sbx;
				end
				6: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h325;
					arA23['h4] = 1'sbx;
				end
				7: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1ed;
					arA23['h4] = 1'sbx;
				end
				8: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1e5;
					arA23['h4] = 1'sbx;
				end
				9: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				10: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				11: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				default: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
			endcase
		else if (opcode[11:6] == 'h23)
			(* full_case, parallel_case *)
			case (col)
				0: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h232;
					arA23['h4] = 1'sbx;
				end
				1: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				2: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h3a0;
					arA23['h4] = 1'sbx;
				end
				3: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				4: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h3a4;
					arA23['h4] = 1'sbx;
				end
				5: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1f1;
					arA23['h4] = 1'sbx;
				end
				6: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h325;
					arA23['h4] = 1'sbx;
				end
				7: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1ed;
					arA23['h4] = 1'sbx;
				end
				8: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1e5;
					arA23['h4] = 1'sbx;
				end
				9: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				10: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				11: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				default: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
			endcase
		else if (opcode[11:6] == 'h28)
			(* full_case, parallel_case *)
			case (col)
				0: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h12d;
					arA23['h4] = 1'sbx;
				end
				1: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				2: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h6;
					arA23['h4] = 'h3c3;
				end
				3: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h21c;
					arA23['h4] = 'h3c3;
				end
				4: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h103;
					arA23['h4] = 'h3c3;
				end
				5: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1c2;
					arA23['h4] = 'h3c3;
				end
				6: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1e3;
					arA23['h4] = 'h3c3;
				end
				7: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'ha;
					arA23['h4] = 'h3c3;
				end
				8: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1e2;
					arA23['h4] = 'h3c3;
				end
				9: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				10: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				11: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				default: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
			endcase
		else if (opcode[11:6] == 'h29)
			(* full_case, parallel_case *)
			case (col)
				0: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h12d;
					arA23['h4] = 1'sbx;
				end
				1: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				2: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h6;
					arA23['h4] = 'h3c3;
				end
				3: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h21c;
					arA23['h4] = 'h3c3;
				end
				4: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h103;
					arA23['h4] = 'h3c3;
				end
				5: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1c2;
					arA23['h4] = 'h3c3;
				end
				6: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1e3;
					arA23['h4] = 'h3c3;
				end
				7: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'ha;
					arA23['h4] = 'h3c3;
				end
				8: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1e2;
					arA23['h4] = 'h3c3;
				end
				9: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				10: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				11: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				default: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
			endcase
		else if (opcode[11:6] == 'h2a)
			(* full_case, parallel_case *)
			case (col)
				0: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h125;
					arA23['h4] = 1'sbx;
				end
				1: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				2: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'hb;
					arA23['h4] = 'h3cb;
				end
				3: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'hf;
					arA23['h4] = 'h3cb;
				end
				4: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h179;
					arA23['h4] = 'h3cb;
				end
				5: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1c6;
					arA23['h4] = 'h3cb;
				end
				6: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1e7;
					arA23['h4] = 'h3cb;
				end
				7: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'he;
					arA23['h4] = 'h3cb;
				end
				8: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1e6;
					arA23['h4] = 'h3cb;
				end
				9: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				10: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				11: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				default: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
			endcase
		else if (opcode[11:6] == 'h2b)
			(* full_case, parallel_case *)
			case (col)
				0: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h345;
					arA23['h4] = 1'sbx;
				end
				1: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				2: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h6;
					arA23['h4] = 'h343;
				end
				3: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h21c;
					arA23['h4] = 'h343;
				end
				4: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h103;
					arA23['h4] = 'h343;
				end
				5: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1c2;
					arA23['h4] = 'h343;
				end
				6: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1e3;
					arA23['h4] = 'h343;
				end
				7: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'ha;
					arA23['h4] = 'h343;
				end
				8: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1e2;
					arA23['h4] = 'h343;
				end
				9: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				10: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				11: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				default: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
			endcase
		else if ((opcode[11:6] & 'h3e) == 'h32)
			(* full_case, parallel_case *)
			case (col)
				0: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				1: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				2: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h127;
					arA23['h4] = 1'sbx;
				end
				3: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h123;
					arA23['h4] = 1'sbx;
				end
				4: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				5: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1fd;
					arA23['h4] = 1'sbx;
				end
				6: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1f5;
					arA23['h4] = 1'sbx;
				end
				7: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1f9;
					arA23['h4] = 1'sbx;
				end
				8: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1e9;
					arA23['h4] = 1'sbx;
				end
				9: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1fd;
					arA23['h4] = 1'sbx;
				end
				10: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1f5;
					arA23['h4] = 1'sbx;
				end
				11: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				default: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
			endcase
		else if ((opcode[11:6] & 'h7) == 'h6)
			(* full_case, parallel_case *)
			case (col)
				0: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h152;
					arA23['h4] = 1'sbx;
				end
				1: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				2: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h6;
					arA23['h4] = 'h151;
				end
				3: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h21c;
					arA23['h4] = 'h151;
				end
				4: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h103;
					arA23['h4] = 'h151;
				end
				5: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1c2;
					arA23['h4] = 'h151;
				end
				6: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1e3;
					arA23['h4] = 'h151;
				end
				7: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'ha;
					arA23['h4] = 'h151;
				end
				8: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1e2;
					arA23['h4] = 'h151;
				end
				9: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1c2;
					arA23['h4] = 'h151;
				end
				10: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1e3;
					arA23['h4] = 'h151;
				end
				11: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'hea;
					arA23['h4] = 'h152;
				end
				default: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
			endcase
		else if ((opcode[11:6] & 'h7) == 'h7)
			(* full_case, parallel_case *)
			case (col)
				0: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				1: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				2: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h2f1;
					arA23['h4] = 1'sbx;
				end
				3: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				4: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				5: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h2f2;
					arA23['h4] = 1'sbx;
				end
				6: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1fb;
					arA23['h4] = 1'sbx;
				end
				7: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h275;
					arA23['h4] = 1'sbx;
				end
				8: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h3e4;
					arA23['h4] = 1'sbx;
				end
				9: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h2f2;
					arA23['h4] = 1'sbx;
				end
				10: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1fb;
					arA23['h4] = 1'sbx;
				end
				11: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				default: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
			endcase
		else if (opcode[11:6] == 'h3a)
			(* full_case, parallel_case *)
			case (col)
				0: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				1: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				2: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h273;
					arA23['h4] = 1'sbx;
				end
				3: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				4: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				5: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h2b0;
					arA23['h4] = 1'sbx;
				end
				6: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1f3;
					arA23['h4] = 1'sbx;
				end
				7: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h293;
					arA23['h4] = 1'sbx;
				end
				8: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1f2;
					arA23['h4] = 1'sbx;
				end
				9: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h2b0;
					arA23['h4] = 1'sbx;
				end
				10: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1f3;
					arA23['h4] = 1'sbx;
				end
				11: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				default: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
			endcase
		else if (opcode[11:6] == 'h3b)
			(* full_case, parallel_case *)
			case (col)
				0: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				1: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				2: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h255;
					arA23['h4] = 1'sbx;
				end
				3: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				4: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				5: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h2b4;
					arA23['h4] = 1'sbx;
				end
				6: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1f7;
					arA23['h4] = 1'sbx;
				end
				7: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h297;
					arA23['h4] = 1'sbx;
				end
				8: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1f6;
					arA23['h4] = 1'sbx;
				end
				9: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h2b4;
					arA23['h4] = 1'sbx;
				end
				10: begin
					arIll['h4] = 1'b0;
					arA1['h4] = 'h1f7;
					arA23['h4] = 1'sbx;
				end
				11: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
				default: begin
					arIll['h4] = 1'b1;
					arA1['h4] = 1'sbx;
					arA23['h4] = 1'sbx;
				end
			endcase
		else if (opcode[11:6] == 'h39) begin
			arIll['h4] = illMisc;
			arA1['h4] = a1Misc;
			arA23['h4] = 1'sbx;
		end
		else begin
			arIll['h4] = 1'b1;
			arA1['h4] = 1'sbx;
			arA23['h4] = 1'sbx;
		end
	end
	always @(*) begin
		if (_sv2v_0)
			;
		(* full_case, parallel_case *)
		case (movEa)
			0:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h121;
						arA23['h1] = 1'sbx;
					end
					1: begin
						arIll['h1] = 1'b1;
						arA1['h1] = 1'sbx;
						arA23['h1] = 1'sbx;
					end
					2: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h6;
						arA23['h1] = 'h29b;
					end
					3: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h21c;
						arA23['h1] = 'h29b;
					end
					4: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h103;
						arA23['h1] = 'h29b;
					end
					5: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h1c2;
						arA23['h1] = 'h29b;
					end
					6: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h1e3;
						arA23['h1] = 'h29b;
					end
					7: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'ha;
						arA23['h1] = 'h29b;
					end
					8: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h1e2;
						arA23['h1] = 'h29b;
					end
					9: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h1c2;
						arA23['h1] = 'h29b;
					end
					10: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h1e3;
						arA23['h1] = 'h29b;
					end
					11: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'hea;
						arA23['h1] = 'h121;
					end
					default: begin
						arIll['h1] = 1'b1;
						arA1['h1] = 1'sbx;
						arA23['h1] = 1'sbx;
					end
				endcase
			2:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h2fa;
						arA23['h1] = 1'sbx;
					end
					1: begin
						arIll['h1] = 1'b1;
						arA1['h1] = 1'sbx;
						arA23['h1] = 1'sbx;
					end
					2: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h6;
						arA23['h1] = 'h3ab;
					end
					3: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h21c;
						arA23['h1] = 'h3ab;
					end
					4: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h103;
						arA23['h1] = 'h3ab;
					end
					5: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h1c2;
						arA23['h1] = 'h3ab;
					end
					6: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h1e3;
						arA23['h1] = 'h3ab;
					end
					7: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'ha;
						arA23['h1] = 'h3ab;
					end
					8: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h1e2;
						arA23['h1] = 'h3ab;
					end
					9: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h1c2;
						arA23['h1] = 'h3ab;
					end
					10: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h1e3;
						arA23['h1] = 'h3ab;
					end
					11: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'hea;
						arA23['h1] = 'h2fa;
					end
					default: begin
						arIll['h1] = 1'b1;
						arA1['h1] = 1'sbx;
						arA23['h1] = 1'sbx;
					end
				endcase
			3:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h2fe;
						arA23['h1] = 1'sbx;
					end
					1: begin
						arIll['h1] = 1'b1;
						arA1['h1] = 1'sbx;
						arA23['h1] = 1'sbx;
					end
					2: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h6;
						arA23['h1] = 'h3af;
					end
					3: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h21c;
						arA23['h1] = 'h3af;
					end
					4: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h103;
						arA23['h1] = 'h3af;
					end
					5: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h1c2;
						arA23['h1] = 'h3af;
					end
					6: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h1e3;
						arA23['h1] = 'h3af;
					end
					7: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'ha;
						arA23['h1] = 'h3af;
					end
					8: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h1e2;
						arA23['h1] = 'h3af;
					end
					9: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h1c2;
						arA23['h1] = 'h3af;
					end
					10: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h1e3;
						arA23['h1] = 'h3af;
					end
					11: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'hea;
						arA23['h1] = 'h2fe;
					end
					default: begin
						arIll['h1] = 1'b1;
						arA1['h1] = 1'sbx;
						arA23['h1] = 1'sbx;
					end
				endcase
			4:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h2f8;
						arA23['h1] = 1'sbx;
					end
					1: begin
						arIll['h1] = 1'b1;
						arA1['h1] = 1'sbx;
						arA23['h1] = 1'sbx;
					end
					2: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h6;
						arA23['h1] = 'h38b;
					end
					3: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h21c;
						arA23['h1] = 'h38b;
					end
					4: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h103;
						arA23['h1] = 'h38b;
					end
					5: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h1c2;
						arA23['h1] = 'h38b;
					end
					6: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h1e3;
						arA23['h1] = 'h38b;
					end
					7: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'ha;
						arA23['h1] = 'h38b;
					end
					8: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h1e2;
						arA23['h1] = 'h38b;
					end
					9: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h1c2;
						arA23['h1] = 'h38b;
					end
					10: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h1e3;
						arA23['h1] = 'h38b;
					end
					11: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'hea;
						arA23['h1] = 'h2f8;
					end
					default: begin
						arIll['h1] = 1'b1;
						arA1['h1] = 1'sbx;
						arA23['h1] = 1'sbx;
					end
				endcase
			5:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h2da;
						arA23['h1] = 1'sbx;
					end
					1: begin
						arIll['h1] = 1'b1;
						arA1['h1] = 1'sbx;
						arA23['h1] = 1'sbx;
					end
					2: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h6;
						arA23['h1] = 'h38a;
					end
					3: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h21c;
						arA23['h1] = 'h38a;
					end
					4: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h103;
						arA23['h1] = 'h38a;
					end
					5: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h1c2;
						arA23['h1] = 'h38a;
					end
					6: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h1e3;
						arA23['h1] = 'h38a;
					end
					7: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'ha;
						arA23['h1] = 'h38a;
					end
					8: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h1e2;
						arA23['h1] = 'h38a;
					end
					9: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h1c2;
						arA23['h1] = 'h38a;
					end
					10: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h1e3;
						arA23['h1] = 'h38a;
					end
					11: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'hea;
						arA23['h1] = 'h2da;
					end
					default: begin
						arIll['h1] = 1'b1;
						arA1['h1] = 1'sbx;
						arA23['h1] = 1'sbx;
					end
				endcase
			6:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h1eb;
						arA23['h1] = 1'sbx;
					end
					1: begin
						arIll['h1] = 1'b1;
						arA1['h1] = 1'sbx;
						arA23['h1] = 1'sbx;
					end
					2: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h6;
						arA23['h1] = 'h298;
					end
					3: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h21c;
						arA23['h1] = 'h298;
					end
					4: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h103;
						arA23['h1] = 'h298;
					end
					5: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h1c2;
						arA23['h1] = 'h298;
					end
					6: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h1e3;
						arA23['h1] = 'h298;
					end
					7: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'ha;
						arA23['h1] = 'h298;
					end
					8: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h1e2;
						arA23['h1] = 'h298;
					end
					9: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h1c2;
						arA23['h1] = 'h298;
					end
					10: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h1e3;
						arA23['h1] = 'h298;
					end
					11: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'hea;
						arA23['h1] = 'h1eb;
					end
					default: begin
						arIll['h1] = 1'b1;
						arA1['h1] = 1'sbx;
						arA23['h1] = 1'sbx;
					end
				endcase
			7:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h2d9;
						arA23['h1] = 1'sbx;
					end
					1: begin
						arIll['h1] = 1'b1;
						arA1['h1] = 1'sbx;
						arA23['h1] = 1'sbx;
					end
					2: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h6;
						arA23['h1] = 'h388;
					end
					3: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h21c;
						arA23['h1] = 'h388;
					end
					4: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h103;
						arA23['h1] = 'h388;
					end
					5: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h1c2;
						arA23['h1] = 'h388;
					end
					6: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h1e3;
						arA23['h1] = 'h388;
					end
					7: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'ha;
						arA23['h1] = 'h388;
					end
					8: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h1e2;
						arA23['h1] = 'h388;
					end
					9: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h1c2;
						arA23['h1] = 'h388;
					end
					10: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h1e3;
						arA23['h1] = 'h388;
					end
					11: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'hea;
						arA23['h1] = 'h2d9;
					end
					default: begin
						arIll['h1] = 1'b1;
						arA1['h1] = 1'sbx;
						arA23['h1] = 1'sbx;
					end
				endcase
			8:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h1ea;
						arA23['h1] = 1'sbx;
					end
					1: begin
						arIll['h1] = 1'b1;
						arA1['h1] = 1'sbx;
						arA23['h1] = 1'sbx;
					end
					2: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h6;
						arA23['h1] = 'h32b;
					end
					3: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h21c;
						arA23['h1] = 'h32b;
					end
					4: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h103;
						arA23['h1] = 'h32b;
					end
					5: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h1c2;
						arA23['h1] = 'h32b;
					end
					6: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h1e3;
						arA23['h1] = 'h32b;
					end
					7: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'ha;
						arA23['h1] = 'h32b;
					end
					8: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h1e2;
						arA23['h1] = 'h32b;
					end
					9: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h1c2;
						arA23['h1] = 'h32b;
					end
					10: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'h1e3;
						arA23['h1] = 'h32b;
					end
					11: begin
						arIll['h1] = 1'b0;
						arA1['h1] = 'hea;
						arA23['h1] = 'h1ea;
					end
					default: begin
						arIll['h1] = 1'b1;
						arA1['h1] = 1'sbx;
						arA23['h1] = 1'sbx;
					end
				endcase
			default: begin
				arIll['h1] = 1'b1;
				arA1['h1] = 1'sbx;
				arA23['h1] = 1'sbx;
			end
		endcase
		(* full_case, parallel_case *)
		case (movEa)
			0:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h129;
						arA23['h2] = 1'sbx;
					end
					1: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h129;
						arA23['h2] = 1'sbx;
					end
					2: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'hb;
						arA23['h2] = 'h29f;
					end
					3: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'hf;
						arA23['h2] = 'h29f;
					end
					4: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h179;
						arA23['h2] = 'h29f;
					end
					5: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h1c6;
						arA23['h2] = 'h29f;
					end
					6: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h1e7;
						arA23['h2] = 'h29f;
					end
					7: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'he;
						arA23['h2] = 'h29f;
					end
					8: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h1e6;
						arA23['h2] = 'h29f;
					end
					9: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h1c6;
						arA23['h2] = 'h29f;
					end
					10: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h1e7;
						arA23['h2] = 'h29f;
					end
					11: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'ha7;
						arA23['h2] = 'h129;
					end
					default: begin
						arIll['h2] = 1'b1;
						arA1['h2] = 1'sbx;
						arA23['h2] = 1'sbx;
					end
				endcase
			1:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h129;
						arA23['h2] = 1'sbx;
					end
					1: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h129;
						arA23['h2] = 1'sbx;
					end
					2: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'hb;
						arA23['h2] = 'h29f;
					end
					3: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'hf;
						arA23['h2] = 'h29f;
					end
					4: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h179;
						arA23['h2] = 'h29f;
					end
					5: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h1c6;
						arA23['h2] = 'h29f;
					end
					6: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h1e7;
						arA23['h2] = 'h29f;
					end
					7: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'he;
						arA23['h2] = 'h29f;
					end
					8: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h1e6;
						arA23['h2] = 'h29f;
					end
					9: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h1c6;
						arA23['h2] = 'h29f;
					end
					10: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h1e7;
						arA23['h2] = 'h29f;
					end
					11: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'ha7;
						arA23['h2] = 'h129;
					end
					default: begin
						arIll['h2] = 1'b1;
						arA1['h2] = 1'sbx;
						arA23['h2] = 1'sbx;
					end
				endcase
			2:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h2f9;
						arA23['h2] = 1'sbx;
					end
					1: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h2f9;
						arA23['h2] = 1'sbx;
					end
					2: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'hb;
						arA23['h2] = 'h3a9;
					end
					3: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'hf;
						arA23['h2] = 'h3a9;
					end
					4: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h179;
						arA23['h2] = 'h3a9;
					end
					5: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h1c6;
						arA23['h2] = 'h3a9;
					end
					6: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h1e7;
						arA23['h2] = 'h3a9;
					end
					7: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'he;
						arA23['h2] = 'h3a9;
					end
					8: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h1e6;
						arA23['h2] = 'h3a9;
					end
					9: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h1c6;
						arA23['h2] = 'h3a9;
					end
					10: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h1e7;
						arA23['h2] = 'h3a9;
					end
					11: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'ha7;
						arA23['h2] = 'h2f9;
					end
					default: begin
						arIll['h2] = 1'b1;
						arA1['h2] = 1'sbx;
						arA23['h2] = 1'sbx;
					end
				endcase
			3:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h2fd;
						arA23['h2] = 1'sbx;
					end
					1: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h2fd;
						arA23['h2] = 1'sbx;
					end
					2: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'hb;
						arA23['h2] = 'h3ad;
					end
					3: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'hf;
						arA23['h2] = 'h3ad;
					end
					4: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h179;
						arA23['h2] = 'h3ad;
					end
					5: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h1c6;
						arA23['h2] = 'h3ad;
					end
					6: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h1e7;
						arA23['h2] = 'h3ad;
					end
					7: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'he;
						arA23['h2] = 'h3ad;
					end
					8: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h1e6;
						arA23['h2] = 'h3ad;
					end
					9: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h1c6;
						arA23['h2] = 'h3ad;
					end
					10: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h1e7;
						arA23['h2] = 'h3ad;
					end
					11: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'ha7;
						arA23['h2] = 'h2fd;
					end
					default: begin
						arIll['h2] = 1'b1;
						arA1['h2] = 1'sbx;
						arA23['h2] = 1'sbx;
					end
				endcase
			4:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h2fc;
						arA23['h2] = 1'sbx;
					end
					1: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h2fc;
						arA23['h2] = 1'sbx;
					end
					2: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'hb;
						arA23['h2] = 'h38f;
					end
					3: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'hf;
						arA23['h2] = 'h38f;
					end
					4: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h179;
						arA23['h2] = 'h38f;
					end
					5: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h1c6;
						arA23['h2] = 'h38f;
					end
					6: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h1e7;
						arA23['h2] = 'h38f;
					end
					7: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'he;
						arA23['h2] = 'h38f;
					end
					8: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h1e6;
						arA23['h2] = 'h38f;
					end
					9: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h1c6;
						arA23['h2] = 'h38f;
					end
					10: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h1e7;
						arA23['h2] = 'h38f;
					end
					11: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'ha7;
						arA23['h2] = 'h2fc;
					end
					default: begin
						arIll['h2] = 1'b1;
						arA1['h2] = 1'sbx;
						arA23['h2] = 1'sbx;
					end
				endcase
			5:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h2de;
						arA23['h2] = 1'sbx;
					end
					1: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h2de;
						arA23['h2] = 1'sbx;
					end
					2: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'hb;
						arA23['h2] = 'h38e;
					end
					3: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'hf;
						arA23['h2] = 'h38e;
					end
					4: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h179;
						arA23['h2] = 'h38e;
					end
					5: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h1c6;
						arA23['h2] = 'h38e;
					end
					6: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h1e7;
						arA23['h2] = 'h38e;
					end
					7: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'he;
						arA23['h2] = 'h38e;
					end
					8: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h1e6;
						arA23['h2] = 'h38e;
					end
					9: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h1c6;
						arA23['h2] = 'h38e;
					end
					10: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h1e7;
						arA23['h2] = 'h38e;
					end
					11: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'ha7;
						arA23['h2] = 'h2de;
					end
					default: begin
						arIll['h2] = 1'b1;
						arA1['h2] = 1'sbx;
						arA23['h2] = 1'sbx;
					end
				endcase
			6:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h1ef;
						arA23['h2] = 1'sbx;
					end
					1: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h1ef;
						arA23['h2] = 1'sbx;
					end
					2: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'hb;
						arA23['h2] = 'h29c;
					end
					3: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'hf;
						arA23['h2] = 'h29c;
					end
					4: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h179;
						arA23['h2] = 'h29c;
					end
					5: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h1c6;
						arA23['h2] = 'h29c;
					end
					6: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h1e7;
						arA23['h2] = 'h29c;
					end
					7: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'he;
						arA23['h2] = 'h29c;
					end
					8: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h1e6;
						arA23['h2] = 'h29c;
					end
					9: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h1c6;
						arA23['h2] = 'h29c;
					end
					10: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h1e7;
						arA23['h2] = 'h29c;
					end
					11: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'ha7;
						arA23['h2] = 'h1ef;
					end
					default: begin
						arIll['h2] = 1'b1;
						arA1['h2] = 1'sbx;
						arA23['h2] = 1'sbx;
					end
				endcase
			7:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h2dd;
						arA23['h2] = 1'sbx;
					end
					1: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h2dd;
						arA23['h2] = 1'sbx;
					end
					2: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'hb;
						arA23['h2] = 'h38c;
					end
					3: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'hf;
						arA23['h2] = 'h38c;
					end
					4: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h179;
						arA23['h2] = 'h38c;
					end
					5: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h1c6;
						arA23['h2] = 'h38c;
					end
					6: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h1e7;
						arA23['h2] = 'h38c;
					end
					7: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'he;
						arA23['h2] = 'h38c;
					end
					8: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h1e6;
						arA23['h2] = 'h38c;
					end
					9: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h1c6;
						arA23['h2] = 'h38c;
					end
					10: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h1e7;
						arA23['h2] = 'h38c;
					end
					11: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'ha7;
						arA23['h2] = 'h2dd;
					end
					default: begin
						arIll['h2] = 1'b1;
						arA1['h2] = 1'sbx;
						arA23['h2] = 1'sbx;
					end
				endcase
			8:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h1ee;
						arA23['h2] = 1'sbx;
					end
					1: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h1ee;
						arA23['h2] = 1'sbx;
					end
					2: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'hb;
						arA23['h2] = 'h30f;
					end
					3: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'hf;
						arA23['h2] = 'h30f;
					end
					4: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h179;
						arA23['h2] = 'h30f;
					end
					5: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h1c6;
						arA23['h2] = 'h30f;
					end
					6: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h1e7;
						arA23['h2] = 'h30f;
					end
					7: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'he;
						arA23['h2] = 'h30f;
					end
					8: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h1e6;
						arA23['h2] = 'h30f;
					end
					9: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h1c6;
						arA23['h2] = 'h30f;
					end
					10: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'h1e7;
						arA23['h2] = 'h30f;
					end
					11: begin
						arIll['h2] = 1'b0;
						arA1['h2] = 'ha7;
						arA23['h2] = 'h1ee;
					end
					default: begin
						arIll['h2] = 1'b1;
						arA1['h2] = 1'sbx;
						arA23['h2] = 1'sbx;
					end
				endcase
			default: begin
				arIll['h2] = 1'b1;
				arA1['h2] = 1'sbx;
				arA23['h2] = 1'sbx;
			end
		endcase
		(* full_case, parallel_case *)
		case (movEa)
			0:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h121;
						arA23['h3] = 1'sbx;
					end
					1: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h121;
						arA23['h3] = 1'sbx;
					end
					2: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h6;
						arA23['h3] = 'h29b;
					end
					3: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h21c;
						arA23['h3] = 'h29b;
					end
					4: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h103;
						arA23['h3] = 'h29b;
					end
					5: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h1c2;
						arA23['h3] = 'h29b;
					end
					6: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h1e3;
						arA23['h3] = 'h29b;
					end
					7: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'ha;
						arA23['h3] = 'h29b;
					end
					8: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h1e2;
						arA23['h3] = 'h29b;
					end
					9: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h1c2;
						arA23['h3] = 'h29b;
					end
					10: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h1e3;
						arA23['h3] = 'h29b;
					end
					11: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'hea;
						arA23['h3] = 'h121;
					end
					default: begin
						arIll['h3] = 1'b1;
						arA1['h3] = 1'sbx;
						arA23['h3] = 1'sbx;
					end
				endcase
			1:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h279;
						arA23['h3] = 1'sbx;
					end
					1: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h279;
						arA23['h3] = 1'sbx;
					end
					2: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h6;
						arA23['h3] = 'h158;
					end
					3: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h21c;
						arA23['h3] = 'h158;
					end
					4: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h103;
						arA23['h3] = 'h158;
					end
					5: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h1c2;
						arA23['h3] = 'h158;
					end
					6: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h1e3;
						arA23['h3] = 'h158;
					end
					7: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'ha;
						arA23['h3] = 'h158;
					end
					8: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h1e2;
						arA23['h3] = 'h158;
					end
					9: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h1c2;
						arA23['h3] = 'h158;
					end
					10: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h1e3;
						arA23['h3] = 'h158;
					end
					11: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'hea;
						arA23['h3] = 'h279;
					end
					default: begin
						arIll['h3] = 1'b1;
						arA1['h3] = 1'sbx;
						arA23['h3] = 1'sbx;
					end
				endcase
			2:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h2fa;
						arA23['h3] = 1'sbx;
					end
					1: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h2fa;
						arA23['h3] = 1'sbx;
					end
					2: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h6;
						arA23['h3] = 'h3ab;
					end
					3: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h21c;
						arA23['h3] = 'h3ab;
					end
					4: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h103;
						arA23['h3] = 'h3ab;
					end
					5: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h1c2;
						arA23['h3] = 'h3ab;
					end
					6: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h1e3;
						arA23['h3] = 'h3ab;
					end
					7: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'ha;
						arA23['h3] = 'h3ab;
					end
					8: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h1e2;
						arA23['h3] = 'h3ab;
					end
					9: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h1c2;
						arA23['h3] = 'h3ab;
					end
					10: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h1e3;
						arA23['h3] = 'h3ab;
					end
					11: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'hea;
						arA23['h3] = 'h2fa;
					end
					default: begin
						arIll['h3] = 1'b1;
						arA1['h3] = 1'sbx;
						arA23['h3] = 1'sbx;
					end
				endcase
			3:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h2fe;
						arA23['h3] = 1'sbx;
					end
					1: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h2fe;
						arA23['h3] = 1'sbx;
					end
					2: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h6;
						arA23['h3] = 'h3af;
					end
					3: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h21c;
						arA23['h3] = 'h3af;
					end
					4: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h103;
						arA23['h3] = 'h3af;
					end
					5: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h1c2;
						arA23['h3] = 'h3af;
					end
					6: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h1e3;
						arA23['h3] = 'h3af;
					end
					7: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'ha;
						arA23['h3] = 'h3af;
					end
					8: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h1e2;
						arA23['h3] = 'h3af;
					end
					9: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h1c2;
						arA23['h3] = 'h3af;
					end
					10: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h1e3;
						arA23['h3] = 'h3af;
					end
					11: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'hea;
						arA23['h3] = 'h2fe;
					end
					default: begin
						arIll['h3] = 1'b1;
						arA1['h3] = 1'sbx;
						arA23['h3] = 1'sbx;
					end
				endcase
			4:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h2f8;
						arA23['h3] = 1'sbx;
					end
					1: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h2f8;
						arA23['h3] = 1'sbx;
					end
					2: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h6;
						arA23['h3] = 'h38b;
					end
					3: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h21c;
						arA23['h3] = 'h38b;
					end
					4: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h103;
						arA23['h3] = 'h38b;
					end
					5: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h1c2;
						arA23['h3] = 'h38b;
					end
					6: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h1e3;
						arA23['h3] = 'h38b;
					end
					7: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'ha;
						arA23['h3] = 'h38b;
					end
					8: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h1e2;
						arA23['h3] = 'h38b;
					end
					9: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h1c2;
						arA23['h3] = 'h38b;
					end
					10: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h1e3;
						arA23['h3] = 'h38b;
					end
					11: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'hea;
						arA23['h3] = 'h2f8;
					end
					default: begin
						arIll['h3] = 1'b1;
						arA1['h3] = 1'sbx;
						arA23['h3] = 1'sbx;
					end
				endcase
			5:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h2da;
						arA23['h3] = 1'sbx;
					end
					1: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h2da;
						arA23['h3] = 1'sbx;
					end
					2: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h6;
						arA23['h3] = 'h38a;
					end
					3: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h21c;
						arA23['h3] = 'h38a;
					end
					4: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h103;
						arA23['h3] = 'h38a;
					end
					5: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h1c2;
						arA23['h3] = 'h38a;
					end
					6: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h1e3;
						arA23['h3] = 'h38a;
					end
					7: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'ha;
						arA23['h3] = 'h38a;
					end
					8: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h1e2;
						arA23['h3] = 'h38a;
					end
					9: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h1c2;
						arA23['h3] = 'h38a;
					end
					10: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h1e3;
						arA23['h3] = 'h38a;
					end
					11: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'hea;
						arA23['h3] = 'h2da;
					end
					default: begin
						arIll['h3] = 1'b1;
						arA1['h3] = 1'sbx;
						arA23['h3] = 1'sbx;
					end
				endcase
			6:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h1eb;
						arA23['h3] = 1'sbx;
					end
					1: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h1eb;
						arA23['h3] = 1'sbx;
					end
					2: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h6;
						arA23['h3] = 'h298;
					end
					3: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h21c;
						arA23['h3] = 'h298;
					end
					4: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h103;
						arA23['h3] = 'h298;
					end
					5: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h1c2;
						arA23['h3] = 'h298;
					end
					6: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h1e3;
						arA23['h3] = 'h298;
					end
					7: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'ha;
						arA23['h3] = 'h298;
					end
					8: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h1e2;
						arA23['h3] = 'h298;
					end
					9: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h1c2;
						arA23['h3] = 'h298;
					end
					10: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h1e3;
						arA23['h3] = 'h298;
					end
					11: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'hea;
						arA23['h3] = 'h1eb;
					end
					default: begin
						arIll['h3] = 1'b1;
						arA1['h3] = 1'sbx;
						arA23['h3] = 1'sbx;
					end
				endcase
			7:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h2d9;
						arA23['h3] = 1'sbx;
					end
					1: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h2d9;
						arA23['h3] = 1'sbx;
					end
					2: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h6;
						arA23['h3] = 'h388;
					end
					3: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h21c;
						arA23['h3] = 'h388;
					end
					4: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h103;
						arA23['h3] = 'h388;
					end
					5: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h1c2;
						arA23['h3] = 'h388;
					end
					6: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h1e3;
						arA23['h3] = 'h388;
					end
					7: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'ha;
						arA23['h3] = 'h388;
					end
					8: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h1e2;
						arA23['h3] = 'h388;
					end
					9: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h1c2;
						arA23['h3] = 'h388;
					end
					10: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h1e3;
						arA23['h3] = 'h388;
					end
					11: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'hea;
						arA23['h3] = 'h2d9;
					end
					default: begin
						arIll['h3] = 1'b1;
						arA1['h3] = 1'sbx;
						arA23['h3] = 1'sbx;
					end
				endcase
			8:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h1ea;
						arA23['h3] = 1'sbx;
					end
					1: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h1ea;
						arA23['h3] = 1'sbx;
					end
					2: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h6;
						arA23['h3] = 'h32b;
					end
					3: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h21c;
						arA23['h3] = 'h32b;
					end
					4: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h103;
						arA23['h3] = 'h32b;
					end
					5: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h1c2;
						arA23['h3] = 'h32b;
					end
					6: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h1e3;
						arA23['h3] = 'h32b;
					end
					7: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'ha;
						arA23['h3] = 'h32b;
					end
					8: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h1e2;
						arA23['h3] = 'h32b;
					end
					9: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h1c2;
						arA23['h3] = 'h32b;
					end
					10: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'h1e3;
						arA23['h3] = 'h32b;
					end
					11: begin
						arIll['h3] = 1'b0;
						arA1['h3] = 'hea;
						arA23['h3] = 'h1ea;
					end
					default: begin
						arIll['h3] = 1'b1;
						arA1['h3] = 1'sbx;
						arA23['h3] = 1'sbx;
					end
				endcase
			default: begin
				arIll['h3] = 1'b1;
				arA1['h3] = 1'sbx;
				arA23['h3] = 1'sbx;
			end
		endcase
		(* full_case, parallel_case *)
		case (row86)
			3'b000:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h2d8;
						arA23['h5] = 1'sbx;
					end
					1: begin
						arIll['h5] = 1'b1;
						arA1['h5] = 1'sbx;
						arA23['h5] = 1'sbx;
					end
					2: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h6;
						arA23['h5] = 'h2f3;
					end
					3: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h21c;
						arA23['h5] = 'h2f3;
					end
					4: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h103;
						arA23['h5] = 'h2f3;
					end
					5: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h1c2;
						arA23['h5] = 'h2f3;
					end
					6: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h1e3;
						arA23['h5] = 'h2f3;
					end
					7: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'ha;
						arA23['h5] = 'h2f3;
					end
					8: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h1e2;
						arA23['h5] = 'h2f3;
					end
					default: begin
						arIll['h5] = 1'b1;
						arA1['h5] = 1'sbx;
						arA23['h5] = 1'sbx;
					end
				endcase
			3'b001:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h2d8;
						arA23['h5] = 1'sbx;
					end
					1: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h2dc;
						arA23['h5] = 1'sbx;
					end
					2: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h6;
						arA23['h5] = 'h2f3;
					end
					3: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h21c;
						arA23['h5] = 'h2f3;
					end
					4: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h103;
						arA23['h5] = 'h2f3;
					end
					5: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h1c2;
						arA23['h5] = 'h2f3;
					end
					6: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h1e3;
						arA23['h5] = 'h2f3;
					end
					7: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'ha;
						arA23['h5] = 'h2f3;
					end
					8: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h1e2;
						arA23['h5] = 'h2f3;
					end
					default: begin
						arIll['h5] = 1'b1;
						arA1['h5] = 1'sbx;
						arA23['h5] = 1'sbx;
					end
				endcase
			3'b010:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h2dc;
						arA23['h5] = 1'sbx;
					end
					1: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h2dc;
						arA23['h5] = 1'sbx;
					end
					2: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'hb;
						arA23['h5] = 'h2f7;
					end
					3: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'hf;
						arA23['h5] = 'h2f7;
					end
					4: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h179;
						arA23['h5] = 'h2f7;
					end
					5: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h1c6;
						arA23['h5] = 'h2f7;
					end
					6: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h1e7;
						arA23['h5] = 'h2f7;
					end
					7: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'he;
						arA23['h5] = 'h2f7;
					end
					8: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h1e6;
						arA23['h5] = 'h2f7;
					end
					default: begin
						arIll['h5] = 1'b1;
						arA1['h5] = 1'sbx;
						arA23['h5] = 1'sbx;
					end
				endcase
			3'b011:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h384;
						arA23['h5] = 1'sbx;
					end
					1: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h6c;
						arA23['h5] = 1'sbx;
					end
					2: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h6;
						arA23['h5] = 'h380;
					end
					3: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h21c;
						arA23['h5] = 'h380;
					end
					4: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h103;
						arA23['h5] = 'h380;
					end
					5: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h1c2;
						arA23['h5] = 'h380;
					end
					6: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h1e3;
						arA23['h5] = 'h380;
					end
					7: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'ha;
						arA23['h5] = 'h380;
					end
					8: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h1e2;
						arA23['h5] = 'h380;
					end
					default: begin
						arIll['h5] = 1'b1;
						arA1['h5] = 1'sbx;
						arA23['h5] = 1'sbx;
					end
				endcase
			3'b100:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h2d8;
						arA23['h5] = 1'sbx;
					end
					1: begin
						arIll['h5] = 1'b1;
						arA1['h5] = 1'sbx;
						arA23['h5] = 1'sbx;
					end
					2: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h6;
						arA23['h5] = 'h2f3;
					end
					3: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h21c;
						arA23['h5] = 'h2f3;
					end
					4: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h103;
						arA23['h5] = 'h2f3;
					end
					5: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h1c2;
						arA23['h5] = 'h2f3;
					end
					6: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h1e3;
						arA23['h5] = 'h2f3;
					end
					7: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'ha;
						arA23['h5] = 'h2f3;
					end
					8: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h1e2;
						arA23['h5] = 'h2f3;
					end
					default: begin
						arIll['h5] = 1'b1;
						arA1['h5] = 1'sbx;
						arA23['h5] = 1'sbx;
					end
				endcase
			3'b101:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h2d8;
						arA23['h5] = 1'sbx;
					end
					1: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h2dc;
						arA23['h5] = 1'sbx;
					end
					2: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h6;
						arA23['h5] = 'h2f3;
					end
					3: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h21c;
						arA23['h5] = 'h2f3;
					end
					4: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h103;
						arA23['h5] = 'h2f3;
					end
					5: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h1c2;
						arA23['h5] = 'h2f3;
					end
					6: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h1e3;
						arA23['h5] = 'h2f3;
					end
					7: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'ha;
						arA23['h5] = 'h2f3;
					end
					8: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h1e2;
						arA23['h5] = 'h2f3;
					end
					default: begin
						arIll['h5] = 1'b1;
						arA1['h5] = 1'sbx;
						arA23['h5] = 1'sbx;
					end
				endcase
			3'b110:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h2dc;
						arA23['h5] = 1'sbx;
					end
					1: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h2dc;
						arA23['h5] = 1'sbx;
					end
					2: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'hb;
						arA23['h5] = 'h2f7;
					end
					3: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'hf;
						arA23['h5] = 'h2f7;
					end
					4: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h179;
						arA23['h5] = 'h2f7;
					end
					5: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h1c6;
						arA23['h5] = 'h2f7;
					end
					6: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h1e7;
						arA23['h5] = 'h2f7;
					end
					7: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'he;
						arA23['h5] = 'h2f7;
					end
					8: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h1e6;
						arA23['h5] = 'h2f7;
					end
					default: begin
						arIll['h5] = 1'b1;
						arA1['h5] = 1'sbx;
						arA23['h5] = 1'sbx;
					end
				endcase
			3'b111:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h384;
						arA23['h5] = 1'sbx;
					end
					1: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h6c;
						arA23['h5] = 1'sbx;
					end
					2: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h6;
						arA23['h5] = 'h380;
					end
					3: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h21c;
						arA23['h5] = 'h380;
					end
					4: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h103;
						arA23['h5] = 'h380;
					end
					5: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h1c2;
						arA23['h5] = 'h380;
					end
					6: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h1e3;
						arA23['h5] = 'h380;
					end
					7: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'ha;
						arA23['h5] = 'h380;
					end
					8: begin
						arIll['h5] = 1'b0;
						arA1['h5] = 'h1e2;
						arA23['h5] = 'h380;
					end
					default: begin
						arIll['h5] = 1'b1;
						arA1['h5] = 1'sbx;
						arA23['h5] = 1'sbx;
					end
				endcase
		endcase
		(* full_case, parallel_case *)
		case (row86)
			3'b000:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h1c1;
						arA23['h8] = 1'sbx;
					end
					1: begin
						arIll['h8] = 1'b1;
						arA1['h8] = 1'sbx;
						arA23['h8] = 1'sbx;
					end
					2: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h6;
						arA23['h8] = 'h1c3;
					end
					3: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h21c;
						arA23['h8] = 'h1c3;
					end
					4: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h103;
						arA23['h8] = 'h1c3;
					end
					5: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h1c2;
						arA23['h8] = 'h1c3;
					end
					6: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h1e3;
						arA23['h8] = 'h1c3;
					end
					7: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'ha;
						arA23['h8] = 'h1c3;
					end
					8: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h1e2;
						arA23['h8] = 'h1c3;
					end
					9: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h1c2;
						arA23['h8] = 'h1c3;
					end
					10: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h1e3;
						arA23['h8] = 'h1c3;
					end
					11: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'hea;
						arA23['h8] = 'h1c1;
					end
					default: begin
						arIll['h8] = 1'b1;
						arA1['h8] = 1'sbx;
						arA23['h8] = 1'sbx;
					end
				endcase
			3'b001:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h1c1;
						arA23['h8] = 1'sbx;
					end
					1: begin
						arIll['h8] = 1'b1;
						arA1['h8] = 1'sbx;
						arA23['h8] = 1'sbx;
					end
					2: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h6;
						arA23['h8] = 'h1c3;
					end
					3: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h21c;
						arA23['h8] = 'h1c3;
					end
					4: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h103;
						arA23['h8] = 'h1c3;
					end
					5: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h1c2;
						arA23['h8] = 'h1c3;
					end
					6: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h1e3;
						arA23['h8] = 'h1c3;
					end
					7: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'ha;
						arA23['h8] = 'h1c3;
					end
					8: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h1e2;
						arA23['h8] = 'h1c3;
					end
					9: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h1c2;
						arA23['h8] = 'h1c3;
					end
					10: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h1e3;
						arA23['h8] = 'h1c3;
					end
					11: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'hea;
						arA23['h8] = 'h1c1;
					end
					default: begin
						arIll['h8] = 1'b1;
						arA1['h8] = 1'sbx;
						arA23['h8] = 1'sbx;
					end
				endcase
			3'b010:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h1c5;
						arA23['h8] = 1'sbx;
					end
					1: begin
						arIll['h8] = 1'b1;
						arA1['h8] = 1'sbx;
						arA23['h8] = 1'sbx;
					end
					2: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'hb;
						arA23['h8] = 'h1cb;
					end
					3: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'hf;
						arA23['h8] = 'h1cb;
					end
					4: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h179;
						arA23['h8] = 'h1cb;
					end
					5: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h1c6;
						arA23['h8] = 'h1cb;
					end
					6: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h1e7;
						arA23['h8] = 'h1cb;
					end
					7: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'he;
						arA23['h8] = 'h1cb;
					end
					8: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h1e6;
						arA23['h8] = 'h1cb;
					end
					9: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h1c6;
						arA23['h8] = 'h1cb;
					end
					10: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h1e7;
						arA23['h8] = 'h1cb;
					end
					11: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'ha7;
						arA23['h8] = 'h1c5;
					end
					default: begin
						arIll['h8] = 1'b1;
						arA1['h8] = 1'sbx;
						arA23['h8] = 1'sbx;
					end
				endcase
			3'b011:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'ha6;
						arA23['h8] = 1'sbx;
					end
					1: begin
						arIll['h8] = 1'b1;
						arA1['h8] = 1'sbx;
						arA23['h8] = 1'sbx;
					end
					2: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h6;
						arA23['h8] = 'ha4;
					end
					3: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h21c;
						arA23['h8] = 'ha4;
					end
					4: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h103;
						arA23['h8] = 'ha4;
					end
					5: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h1c2;
						arA23['h8] = 'ha4;
					end
					6: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h1e3;
						arA23['h8] = 'ha4;
					end
					7: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'ha;
						arA23['h8] = 'ha4;
					end
					8: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h1e2;
						arA23['h8] = 'ha4;
					end
					9: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h1c2;
						arA23['h8] = 'ha4;
					end
					10: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h1e3;
						arA23['h8] = 'ha4;
					end
					11: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'hea;
						arA23['h8] = 'ha6;
					end
					default: begin
						arIll['h8] = 1'b1;
						arA1['h8] = 1'sbx;
						arA23['h8] = 1'sbx;
					end
				endcase
			3'b100:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h1cd;
						arA23['h8] = 1'sbx;
					end
					1: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h107;
						arA23['h8] = 1'sbx;
					end
					2: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h6;
						arA23['h8] = 'h299;
					end
					3: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h21c;
						arA23['h8] = 'h299;
					end
					4: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h103;
						arA23['h8] = 'h299;
					end
					5: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h1c2;
						arA23['h8] = 'h299;
					end
					6: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h1e3;
						arA23['h8] = 'h299;
					end
					7: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'ha;
						arA23['h8] = 'h299;
					end
					8: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h1e2;
						arA23['h8] = 'h299;
					end
					9: begin
						arIll['h8] = 1'b1;
						arA1['h8] = 1'sbx;
						arA23['h8] = 1'sbx;
					end
					10: begin
						arIll['h8] = 1'b1;
						arA1['h8] = 1'sbx;
						arA23['h8] = 1'sbx;
					end
					11: begin
						arIll['h8] = 1'b1;
						arA1['h8] = 1'sbx;
						arA23['h8] = 1'sbx;
					end
					default: begin
						arIll['h8] = 1'b1;
						arA1['h8] = 1'sbx;
						arA23['h8] = 1'sbx;
					end
				endcase
			3'b101:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['h8] = 1'b1;
						arA1['h8] = 1'sbx;
						arA23['h8] = 1'sbx;
					end
					1: begin
						arIll['h8] = 1'b1;
						arA1['h8] = 1'sbx;
						arA23['h8] = 1'sbx;
					end
					2: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h6;
						arA23['h8] = 'h299;
					end
					3: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h21c;
						arA23['h8] = 'h299;
					end
					4: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h103;
						arA23['h8] = 'h299;
					end
					5: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h1c2;
						arA23['h8] = 'h299;
					end
					6: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h1e3;
						arA23['h8] = 'h299;
					end
					7: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'ha;
						arA23['h8] = 'h299;
					end
					8: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h1e2;
						arA23['h8] = 'h299;
					end
					9: begin
						arIll['h8] = 1'b1;
						arA1['h8] = 1'sbx;
						arA23['h8] = 1'sbx;
					end
					10: begin
						arIll['h8] = 1'b1;
						arA1['h8] = 1'sbx;
						arA23['h8] = 1'sbx;
					end
					11: begin
						arIll['h8] = 1'b1;
						arA1['h8] = 1'sbx;
						arA23['h8] = 1'sbx;
					end
					default: begin
						arIll['h8] = 1'b1;
						arA1['h8] = 1'sbx;
						arA23['h8] = 1'sbx;
					end
				endcase
			3'b110:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['h8] = 1'b1;
						arA1['h8] = 1'sbx;
						arA23['h8] = 1'sbx;
					end
					1: begin
						arIll['h8] = 1'b1;
						arA1['h8] = 1'sbx;
						arA23['h8] = 1'sbx;
					end
					2: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'hb;
						arA23['h8] = 'h29d;
					end
					3: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'hf;
						arA23['h8] = 'h29d;
					end
					4: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h179;
						arA23['h8] = 'h29d;
					end
					5: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h1c6;
						arA23['h8] = 'h29d;
					end
					6: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h1e7;
						arA23['h8] = 'h29d;
					end
					7: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'he;
						arA23['h8] = 'h29d;
					end
					8: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h1e6;
						arA23['h8] = 'h29d;
					end
					9: begin
						arIll['h8] = 1'b1;
						arA1['h8] = 1'sbx;
						arA23['h8] = 1'sbx;
					end
					10: begin
						arIll['h8] = 1'b1;
						arA1['h8] = 1'sbx;
						arA23['h8] = 1'sbx;
					end
					11: begin
						arIll['h8] = 1'b1;
						arA1['h8] = 1'sbx;
						arA23['h8] = 1'sbx;
					end
					default: begin
						arIll['h8] = 1'b1;
						arA1['h8] = 1'sbx;
						arA23['h8] = 1'sbx;
					end
				endcase
			3'b111:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'hae;
						arA23['h8] = 1'sbx;
					end
					1: begin
						arIll['h8] = 1'b1;
						arA1['h8] = 1'sbx;
						arA23['h8] = 1'sbx;
					end
					2: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h6;
						arA23['h8] = 'hac;
					end
					3: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h21c;
						arA23['h8] = 'hac;
					end
					4: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h103;
						arA23['h8] = 'hac;
					end
					5: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h1c2;
						arA23['h8] = 'hac;
					end
					6: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h1e3;
						arA23['h8] = 'hac;
					end
					7: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'ha;
						arA23['h8] = 'hac;
					end
					8: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h1e2;
						arA23['h8] = 'hac;
					end
					9: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h1c2;
						arA23['h8] = 'hac;
					end
					10: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'h1e3;
						arA23['h8] = 'hac;
					end
					11: begin
						arIll['h8] = 1'b0;
						arA1['h8] = 'hea;
						arA23['h8] = 'hae;
					end
					default: begin
						arIll['h8] = 1'b1;
						arA1['h8] = 1'sbx;
						arA23['h8] = 1'sbx;
					end
				endcase
		endcase
		(* full_case, parallel_case *)
		case (row86)
			3'b000:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h1c1;
						arA23['h9] = 1'sbx;
					end
					1: begin
						arIll['h9] = 1'b1;
						arA1['h9] = 1'sbx;
						arA23['h9] = 1'sbx;
					end
					2: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h6;
						arA23['h9] = 'h1c3;
					end
					3: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h21c;
						arA23['h9] = 'h1c3;
					end
					4: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h103;
						arA23['h9] = 'h1c3;
					end
					5: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h1c2;
						arA23['h9] = 'h1c3;
					end
					6: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h1e3;
						arA23['h9] = 'h1c3;
					end
					7: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'ha;
						arA23['h9] = 'h1c3;
					end
					8: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h1e2;
						arA23['h9] = 'h1c3;
					end
					9: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h1c2;
						arA23['h9] = 'h1c3;
					end
					10: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h1e3;
						arA23['h9] = 'h1c3;
					end
					11: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'hea;
						arA23['h9] = 'h1c1;
					end
					default: begin
						arIll['h9] = 1'b1;
						arA1['h9] = 1'sbx;
						arA23['h9] = 1'sbx;
					end
				endcase
			3'b001:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h1c1;
						arA23['h9] = 1'sbx;
					end
					1: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h1c1;
						arA23['h9] = 1'sbx;
					end
					2: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h6;
						arA23['h9] = 'h1c3;
					end
					3: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h21c;
						arA23['h9] = 'h1c3;
					end
					4: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h103;
						arA23['h9] = 'h1c3;
					end
					5: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h1c2;
						arA23['h9] = 'h1c3;
					end
					6: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h1e3;
						arA23['h9] = 'h1c3;
					end
					7: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'ha;
						arA23['h9] = 'h1c3;
					end
					8: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h1e2;
						arA23['h9] = 'h1c3;
					end
					9: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h1c2;
						arA23['h9] = 'h1c3;
					end
					10: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h1e3;
						arA23['h9] = 'h1c3;
					end
					11: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'hea;
						arA23['h9] = 'h1c1;
					end
					default: begin
						arIll['h9] = 1'b1;
						arA1['h9] = 1'sbx;
						arA23['h9] = 1'sbx;
					end
				endcase
			3'b010:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h1c5;
						arA23['h9] = 1'sbx;
					end
					1: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h1c5;
						arA23['h9] = 1'sbx;
					end
					2: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'hb;
						arA23['h9] = 'h1cb;
					end
					3: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'hf;
						arA23['h9] = 'h1cb;
					end
					4: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h179;
						arA23['h9] = 'h1cb;
					end
					5: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h1c6;
						arA23['h9] = 'h1cb;
					end
					6: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h1e7;
						arA23['h9] = 'h1cb;
					end
					7: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'he;
						arA23['h9] = 'h1cb;
					end
					8: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h1e6;
						arA23['h9] = 'h1cb;
					end
					9: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h1c6;
						arA23['h9] = 'h1cb;
					end
					10: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h1e7;
						arA23['h9] = 'h1cb;
					end
					11: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'ha7;
						arA23['h9] = 'h1c5;
					end
					default: begin
						arIll['h9] = 1'b1;
						arA1['h9] = 1'sbx;
						arA23['h9] = 1'sbx;
					end
				endcase
			3'b011:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h1c9;
						arA23['h9] = 1'sbx;
					end
					1: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h1c9;
						arA23['h9] = 1'sbx;
					end
					2: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h6;
						arA23['h9] = 'h1c7;
					end
					3: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h21c;
						arA23['h9] = 'h1c7;
					end
					4: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h103;
						arA23['h9] = 'h1c7;
					end
					5: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h1c2;
						arA23['h9] = 'h1c7;
					end
					6: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h1e3;
						arA23['h9] = 'h1c7;
					end
					7: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'ha;
						arA23['h9] = 'h1c7;
					end
					8: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h1e2;
						arA23['h9] = 'h1c7;
					end
					9: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h1c2;
						arA23['h9] = 'h1c7;
					end
					10: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h1e3;
						arA23['h9] = 'h1c7;
					end
					11: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'hea;
						arA23['h9] = 'h1c9;
					end
					default: begin
						arIll['h9] = 1'b1;
						arA1['h9] = 1'sbx;
						arA23['h9] = 1'sbx;
					end
				endcase
			3'b100:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h1c1;
						arA23['h9] = 1'sbx;
					end
					1: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h10f;
						arA23['h9] = 1'sbx;
					end
					2: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h6;
						arA23['h9] = 'h299;
					end
					3: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h21c;
						arA23['h9] = 'h299;
					end
					4: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h103;
						arA23['h9] = 'h299;
					end
					5: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h1c2;
						arA23['h9] = 'h299;
					end
					6: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h1e3;
						arA23['h9] = 'h299;
					end
					7: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'ha;
						arA23['h9] = 'h299;
					end
					8: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h1e2;
						arA23['h9] = 'h299;
					end
					9: begin
						arIll['h9] = 1'b1;
						arA1['h9] = 1'sbx;
						arA23['h9] = 1'sbx;
					end
					10: begin
						arIll['h9] = 1'b1;
						arA1['h9] = 1'sbx;
						arA23['h9] = 1'sbx;
					end
					11: begin
						arIll['h9] = 1'b1;
						arA1['h9] = 1'sbx;
						arA23['h9] = 1'sbx;
					end
					default: begin
						arIll['h9] = 1'b1;
						arA1['h9] = 1'sbx;
						arA23['h9] = 1'sbx;
					end
				endcase
			3'b101:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h1c1;
						arA23['h9] = 1'sbx;
					end
					1: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h10f;
						arA23['h9] = 1'sbx;
					end
					2: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h6;
						arA23['h9] = 'h299;
					end
					3: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h21c;
						arA23['h9] = 'h299;
					end
					4: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h103;
						arA23['h9] = 'h299;
					end
					5: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h1c2;
						arA23['h9] = 'h299;
					end
					6: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h1e3;
						arA23['h9] = 'h299;
					end
					7: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'ha;
						arA23['h9] = 'h299;
					end
					8: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h1e2;
						arA23['h9] = 'h299;
					end
					9: begin
						arIll['h9] = 1'b1;
						arA1['h9] = 1'sbx;
						arA23['h9] = 1'sbx;
					end
					10: begin
						arIll['h9] = 1'b1;
						arA1['h9] = 1'sbx;
						arA23['h9] = 1'sbx;
					end
					11: begin
						arIll['h9] = 1'b1;
						arA1['h9] = 1'sbx;
						arA23['h9] = 1'sbx;
					end
					default: begin
						arIll['h9] = 1'b1;
						arA1['h9] = 1'sbx;
						arA23['h9] = 1'sbx;
					end
				endcase
			3'b110:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h1c5;
						arA23['h9] = 1'sbx;
					end
					1: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h10b;
						arA23['h9] = 1'sbx;
					end
					2: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'hb;
						arA23['h9] = 'h29d;
					end
					3: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'hf;
						arA23['h9] = 'h29d;
					end
					4: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h179;
						arA23['h9] = 'h29d;
					end
					5: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h1c6;
						arA23['h9] = 'h29d;
					end
					6: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h1e7;
						arA23['h9] = 'h29d;
					end
					7: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'he;
						arA23['h9] = 'h29d;
					end
					8: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h1e6;
						arA23['h9] = 'h29d;
					end
					9: begin
						arIll['h9] = 1'b1;
						arA1['h9] = 1'sbx;
						arA23['h9] = 1'sbx;
					end
					10: begin
						arIll['h9] = 1'b1;
						arA1['h9] = 1'sbx;
						arA23['h9] = 1'sbx;
					end
					11: begin
						arIll['h9] = 1'b1;
						arA1['h9] = 1'sbx;
						arA23['h9] = 1'sbx;
					end
					default: begin
						arIll['h9] = 1'b1;
						arA1['h9] = 1'sbx;
						arA23['h9] = 1'sbx;
					end
				endcase
			3'b111:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h1c5;
						arA23['h9] = 1'sbx;
					end
					1: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h1c5;
						arA23['h9] = 1'sbx;
					end
					2: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'hb;
						arA23['h9] = 'h1cb;
					end
					3: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'hf;
						arA23['h9] = 'h1cb;
					end
					4: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h179;
						arA23['h9] = 'h1cb;
					end
					5: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h1c6;
						arA23['h9] = 'h1cb;
					end
					6: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h1e7;
						arA23['h9] = 'h1cb;
					end
					7: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'he;
						arA23['h9] = 'h1cb;
					end
					8: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h1e6;
						arA23['h9] = 'h1cb;
					end
					9: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h1c6;
						arA23['h9] = 'h1cb;
					end
					10: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'h1e7;
						arA23['h9] = 'h1cb;
					end
					11: begin
						arIll['h9] = 1'b0;
						arA1['h9] = 'ha7;
						arA23['h9] = 'h1c5;
					end
					default: begin
						arIll['h9] = 1'b1;
						arA1['h9] = 1'sbx;
						arA23['h9] = 1'sbx;
					end
				endcase
		endcase
		(* full_case, parallel_case *)
		case (row86)
			3'b000:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h1d1;
						arA23['hb] = 1'sbx;
					end
					1: begin
						arIll['hb] = 1'b1;
						arA1['hb] = 1'sbx;
						arA23['hb] = 1'sbx;
					end
					2: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h6;
						arA23['hb] = 'h1d3;
					end
					3: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h21c;
						arA23['hb] = 'h1d3;
					end
					4: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h103;
						arA23['hb] = 'h1d3;
					end
					5: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h1c2;
						arA23['hb] = 'h1d3;
					end
					6: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h1e3;
						arA23['hb] = 'h1d3;
					end
					7: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'ha;
						arA23['hb] = 'h1d3;
					end
					8: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h1e2;
						arA23['hb] = 'h1d3;
					end
					9: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h1c2;
						arA23['hb] = 'h1d3;
					end
					10: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h1e3;
						arA23['hb] = 'h1d3;
					end
					11: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'hea;
						arA23['hb] = 'h1d1;
					end
					default: begin
						arIll['hb] = 1'b1;
						arA1['hb] = 1'sbx;
						arA23['hb] = 1'sbx;
					end
				endcase
			3'b001:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h1d1;
						arA23['hb] = 1'sbx;
					end
					1: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h1d1;
						arA23['hb] = 1'sbx;
					end
					2: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h6;
						arA23['hb] = 'h1d3;
					end
					3: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h21c;
						arA23['hb] = 'h1d3;
					end
					4: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h103;
						arA23['hb] = 'h1d3;
					end
					5: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h1c2;
						arA23['hb] = 'h1d3;
					end
					6: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h1e3;
						arA23['hb] = 'h1d3;
					end
					7: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'ha;
						arA23['hb] = 'h1d3;
					end
					8: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h1e2;
						arA23['hb] = 'h1d3;
					end
					9: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h1c2;
						arA23['hb] = 'h1d3;
					end
					10: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h1e3;
						arA23['hb] = 'h1d3;
					end
					11: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'hea;
						arA23['hb] = 'h1d1;
					end
					default: begin
						arIll['hb] = 1'b1;
						arA1['hb] = 1'sbx;
						arA23['hb] = 1'sbx;
					end
				endcase
			3'b010:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h1d5;
						arA23['hb] = 1'sbx;
					end
					1: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h1d5;
						arA23['hb] = 1'sbx;
					end
					2: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'hb;
						arA23['hb] = 'h1d7;
					end
					3: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'hf;
						arA23['hb] = 'h1d7;
					end
					4: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h179;
						arA23['hb] = 'h1d7;
					end
					5: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h1c6;
						arA23['hb] = 'h1d7;
					end
					6: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h1e7;
						arA23['hb] = 'h1d7;
					end
					7: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'he;
						arA23['hb] = 'h1d7;
					end
					8: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h1e6;
						arA23['hb] = 'h1d7;
					end
					9: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h1c6;
						arA23['hb] = 'h1d7;
					end
					10: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h1e7;
						arA23['hb] = 'h1d7;
					end
					11: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'ha7;
						arA23['hb] = 'h1d5;
					end
					default: begin
						arIll['hb] = 1'b1;
						arA1['hb] = 1'sbx;
						arA23['hb] = 1'sbx;
					end
				endcase
			3'b011:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h1d9;
						arA23['hb] = 1'sbx;
					end
					1: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h1d9;
						arA23['hb] = 1'sbx;
					end
					2: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h6;
						arA23['hb] = 'h1cf;
					end
					3: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h21c;
						arA23['hb] = 'h1cf;
					end
					4: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h103;
						arA23['hb] = 'h1cf;
					end
					5: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h1c2;
						arA23['hb] = 'h1cf;
					end
					6: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h1e3;
						arA23['hb] = 'h1cf;
					end
					7: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'ha;
						arA23['hb] = 'h1cf;
					end
					8: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h1e2;
						arA23['hb] = 'h1cf;
					end
					9: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h1c2;
						arA23['hb] = 'h1cf;
					end
					10: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h1e3;
						arA23['hb] = 'h1cf;
					end
					11: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'hea;
						arA23['hb] = 'h1d9;
					end
					default: begin
						arIll['hb] = 1'b1;
						arA1['hb] = 1'sbx;
						arA23['hb] = 1'sbx;
					end
				endcase
			3'b100:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h100;
						arA23['hb] = 1'sbx;
					end
					1: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h6b;
						arA23['hb] = 1'sbx;
					end
					2: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h6;
						arA23['hb] = 'h299;
					end
					3: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h21c;
						arA23['hb] = 'h299;
					end
					4: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h103;
						arA23['hb] = 'h299;
					end
					5: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h1c2;
						arA23['hb] = 'h299;
					end
					6: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h1e3;
						arA23['hb] = 'h299;
					end
					7: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'ha;
						arA23['hb] = 'h299;
					end
					8: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h1e2;
						arA23['hb] = 'h299;
					end
					9: begin
						arIll['hb] = 1'b1;
						arA1['hb] = 1'sbx;
						arA23['hb] = 1'sbx;
					end
					10: begin
						arIll['hb] = 1'b1;
						arA1['hb] = 1'sbx;
						arA23['hb] = 1'sbx;
					end
					11: begin
						arIll['hb] = 1'b1;
						arA1['hb] = 1'sbx;
						arA23['hb] = 1'sbx;
					end
					default: begin
						arIll['hb] = 1'b1;
						arA1['hb] = 1'sbx;
						arA23['hb] = 1'sbx;
					end
				endcase
			3'b101:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h100;
						arA23['hb] = 1'sbx;
					end
					1: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h6b;
						arA23['hb] = 1'sbx;
					end
					2: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h6;
						arA23['hb] = 'h299;
					end
					3: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h21c;
						arA23['hb] = 'h299;
					end
					4: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h103;
						arA23['hb] = 'h299;
					end
					5: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h1c2;
						arA23['hb] = 'h299;
					end
					6: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h1e3;
						arA23['hb] = 'h299;
					end
					7: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'ha;
						arA23['hb] = 'h299;
					end
					8: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h1e2;
						arA23['hb] = 'h299;
					end
					9: begin
						arIll['hb] = 1'b1;
						arA1['hb] = 1'sbx;
						arA23['hb] = 1'sbx;
					end
					10: begin
						arIll['hb] = 1'b1;
						arA1['hb] = 1'sbx;
						arA23['hb] = 1'sbx;
					end
					11: begin
						arIll['hb] = 1'b1;
						arA1['hb] = 1'sbx;
						arA23['hb] = 1'sbx;
					end
					default: begin
						arIll['hb] = 1'b1;
						arA1['hb] = 1'sbx;
						arA23['hb] = 1'sbx;
					end
				endcase
			3'b110:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h10c;
						arA23['hb] = 1'sbx;
					end
					1: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h6f;
						arA23['hb] = 1'sbx;
					end
					2: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'hb;
						arA23['hb] = 'h29d;
					end
					3: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'hf;
						arA23['hb] = 'h29d;
					end
					4: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h179;
						arA23['hb] = 'h29d;
					end
					5: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h1c6;
						arA23['hb] = 'h29d;
					end
					6: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h1e7;
						arA23['hb] = 'h29d;
					end
					7: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'he;
						arA23['hb] = 'h29d;
					end
					8: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h1e6;
						arA23['hb] = 'h29d;
					end
					9: begin
						arIll['hb] = 1'b1;
						arA1['hb] = 1'sbx;
						arA23['hb] = 1'sbx;
					end
					10: begin
						arIll['hb] = 1'b1;
						arA1['hb] = 1'sbx;
						arA23['hb] = 1'sbx;
					end
					11: begin
						arIll['hb] = 1'b1;
						arA1['hb] = 1'sbx;
						arA23['hb] = 1'sbx;
					end
					default: begin
						arIll['hb] = 1'b1;
						arA1['hb] = 1'sbx;
						arA23['hb] = 1'sbx;
					end
				endcase
			3'b111:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h1d5;
						arA23['hb] = 1'sbx;
					end
					1: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h1d5;
						arA23['hb] = 1'sbx;
					end
					2: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'hb;
						arA23['hb] = 'h1d7;
					end
					3: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'hf;
						arA23['hb] = 'h1d7;
					end
					4: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h179;
						arA23['hb] = 'h1d7;
					end
					5: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h1c6;
						arA23['hb] = 'h1d7;
					end
					6: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h1e7;
						arA23['hb] = 'h1d7;
					end
					7: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'he;
						arA23['hb] = 'h1d7;
					end
					8: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h1e6;
						arA23['hb] = 'h1d7;
					end
					9: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h1c6;
						arA23['hb] = 'h1d7;
					end
					10: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'h1e7;
						arA23['hb] = 'h1d7;
					end
					11: begin
						arIll['hb] = 1'b0;
						arA1['hb] = 'ha7;
						arA23['hb] = 'h1d5;
					end
					default: begin
						arIll['hb] = 1'b1;
						arA1['hb] = 1'sbx;
						arA23['hb] = 1'sbx;
					end
				endcase
		endcase
		(* full_case, parallel_case *)
		case (row86)
			3'b000:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h1c1;
						arA23['hc] = 1'sbx;
					end
					1: begin
						arIll['hc] = 1'b1;
						arA1['hc] = 1'sbx;
						arA23['hc] = 1'sbx;
					end
					2: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h6;
						arA23['hc] = 'h1c3;
					end
					3: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h21c;
						arA23['hc] = 'h1c3;
					end
					4: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h103;
						arA23['hc] = 'h1c3;
					end
					5: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h1c2;
						arA23['hc] = 'h1c3;
					end
					6: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h1e3;
						arA23['hc] = 'h1c3;
					end
					7: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'ha;
						arA23['hc] = 'h1c3;
					end
					8: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h1e2;
						arA23['hc] = 'h1c3;
					end
					9: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h1c2;
						arA23['hc] = 'h1c3;
					end
					10: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h1e3;
						arA23['hc] = 'h1c3;
					end
					11: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'hea;
						arA23['hc] = 'h1c1;
					end
					default: begin
						arIll['hc] = 1'b1;
						arA1['hc] = 1'sbx;
						arA23['hc] = 1'sbx;
					end
				endcase
			3'b001:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h1c1;
						arA23['hc] = 1'sbx;
					end
					1: begin
						arIll['hc] = 1'b1;
						arA1['hc] = 1'sbx;
						arA23['hc] = 1'sbx;
					end
					2: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h6;
						arA23['hc] = 'h1c3;
					end
					3: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h21c;
						arA23['hc] = 'h1c3;
					end
					4: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h103;
						arA23['hc] = 'h1c3;
					end
					5: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h1c2;
						arA23['hc] = 'h1c3;
					end
					6: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h1e3;
						arA23['hc] = 'h1c3;
					end
					7: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'ha;
						arA23['hc] = 'h1c3;
					end
					8: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h1e2;
						arA23['hc] = 'h1c3;
					end
					9: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h1c2;
						arA23['hc] = 'h1c3;
					end
					10: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h1e3;
						arA23['hc] = 'h1c3;
					end
					11: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'hea;
						arA23['hc] = 'h1c1;
					end
					default: begin
						arIll['hc] = 1'b1;
						arA1['hc] = 1'sbx;
						arA23['hc] = 1'sbx;
					end
				endcase
			3'b010:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h1c5;
						arA23['hc] = 1'sbx;
					end
					1: begin
						arIll['hc] = 1'b1;
						arA1['hc] = 1'sbx;
						arA23['hc] = 1'sbx;
					end
					2: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'hb;
						arA23['hc] = 'h1cb;
					end
					3: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'hf;
						arA23['hc] = 'h1cb;
					end
					4: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h179;
						arA23['hc] = 'h1cb;
					end
					5: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h1c6;
						arA23['hc] = 'h1cb;
					end
					6: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h1e7;
						arA23['hc] = 'h1cb;
					end
					7: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'he;
						arA23['hc] = 'h1cb;
					end
					8: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h1e6;
						arA23['hc] = 'h1cb;
					end
					9: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h1c6;
						arA23['hc] = 'h1cb;
					end
					10: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h1e7;
						arA23['hc] = 'h1cb;
					end
					11: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'ha7;
						arA23['hc] = 'h1c5;
					end
					default: begin
						arIll['hc] = 1'b1;
						arA1['hc] = 1'sbx;
						arA23['hc] = 1'sbx;
					end
				endcase
			3'b011:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h15b;
						arA23['hc] = 1'sbx;
					end
					1: begin
						arIll['hc] = 1'b1;
						arA1['hc] = 1'sbx;
						arA23['hc] = 1'sbx;
					end
					2: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h6;
						arA23['hc] = 'h15a;
					end
					3: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h21c;
						arA23['hc] = 'h15a;
					end
					4: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h103;
						arA23['hc] = 'h15a;
					end
					5: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h1c2;
						arA23['hc] = 'h15a;
					end
					6: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h1e3;
						arA23['hc] = 'h15a;
					end
					7: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'ha;
						arA23['hc] = 'h15a;
					end
					8: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h1e2;
						arA23['hc] = 'h15a;
					end
					9: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h1c2;
						arA23['hc] = 'h15a;
					end
					10: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h1e3;
						arA23['hc] = 'h15a;
					end
					11: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'hea;
						arA23['hc] = 'h15b;
					end
					default: begin
						arIll['hc] = 1'b1;
						arA1['hc] = 1'sbx;
						arA23['hc] = 1'sbx;
					end
				endcase
			3'b100:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h1cd;
						arA23['hc] = 1'sbx;
					end
					1: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h107;
						arA23['hc] = 1'sbx;
					end
					2: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h6;
						arA23['hc] = 'h299;
					end
					3: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h21c;
						arA23['hc] = 'h299;
					end
					4: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h103;
						arA23['hc] = 'h299;
					end
					5: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h1c2;
						arA23['hc] = 'h299;
					end
					6: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h1e3;
						arA23['hc] = 'h299;
					end
					7: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'ha;
						arA23['hc] = 'h299;
					end
					8: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h1e2;
						arA23['hc] = 'h299;
					end
					9: begin
						arIll['hc] = 1'b1;
						arA1['hc] = 1'sbx;
						arA23['hc] = 1'sbx;
					end
					10: begin
						arIll['hc] = 1'b1;
						arA1['hc] = 1'sbx;
						arA23['hc] = 1'sbx;
					end
					11: begin
						arIll['hc] = 1'b1;
						arA1['hc] = 1'sbx;
						arA23['hc] = 1'sbx;
					end
					default: begin
						arIll['hc] = 1'b1;
						arA1['hc] = 1'sbx;
						arA23['hc] = 1'sbx;
					end
				endcase
			3'b101:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h3e3;
						arA23['hc] = 1'sbx;
					end
					1: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h3e3;
						arA23['hc] = 1'sbx;
					end
					2: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h6;
						arA23['hc] = 'h299;
					end
					3: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h21c;
						arA23['hc] = 'h299;
					end
					4: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h103;
						arA23['hc] = 'h299;
					end
					5: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h1c2;
						arA23['hc] = 'h299;
					end
					6: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h1e3;
						arA23['hc] = 'h299;
					end
					7: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'ha;
						arA23['hc] = 'h299;
					end
					8: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h1e2;
						arA23['hc] = 'h299;
					end
					9: begin
						arIll['hc] = 1'b1;
						arA1['hc] = 1'sbx;
						arA23['hc] = 1'sbx;
					end
					10: begin
						arIll['hc] = 1'b1;
						arA1['hc] = 1'sbx;
						arA23['hc] = 1'sbx;
					end
					11: begin
						arIll['hc] = 1'b1;
						arA1['hc] = 1'sbx;
						arA23['hc] = 1'sbx;
					end
					default: begin
						arIll['hc] = 1'b1;
						arA1['hc] = 1'sbx;
						arA23['hc] = 1'sbx;
					end
				endcase
			3'b110:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['hc] = 1'b1;
						arA1['hc] = 1'sbx;
						arA23['hc] = 1'sbx;
					end
					1: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h3e3;
						arA23['hc] = 1'sbx;
					end
					2: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'hb;
						arA23['hc] = 'h29d;
					end
					3: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'hf;
						arA23['hc] = 'h29d;
					end
					4: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h179;
						arA23['hc] = 'h29d;
					end
					5: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h1c6;
						arA23['hc] = 'h29d;
					end
					6: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h1e7;
						arA23['hc] = 'h29d;
					end
					7: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'he;
						arA23['hc] = 'h29d;
					end
					8: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h1e6;
						arA23['hc] = 'h29d;
					end
					9: begin
						arIll['hc] = 1'b1;
						arA1['hc] = 1'sbx;
						arA23['hc] = 1'sbx;
					end
					10: begin
						arIll['hc] = 1'b1;
						arA1['hc] = 1'sbx;
						arA23['hc] = 1'sbx;
					end
					11: begin
						arIll['hc] = 1'b1;
						arA1['hc] = 1'sbx;
						arA23['hc] = 1'sbx;
					end
					default: begin
						arIll['hc] = 1'b1;
						arA1['hc] = 1'sbx;
						arA23['hc] = 1'sbx;
					end
				endcase
			3'b111:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h15b;
						arA23['hc] = 1'sbx;
					end
					1: begin
						arIll['hc] = 1'b1;
						arA1['hc] = 1'sbx;
						arA23['hc] = 1'sbx;
					end
					2: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h6;
						arA23['hc] = 'h15a;
					end
					3: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h21c;
						arA23['hc] = 'h15a;
					end
					4: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h103;
						arA23['hc] = 'h15a;
					end
					5: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h1c2;
						arA23['hc] = 'h15a;
					end
					6: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h1e3;
						arA23['hc] = 'h15a;
					end
					7: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'ha;
						arA23['hc] = 'h15a;
					end
					8: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h1e2;
						arA23['hc] = 'h15a;
					end
					9: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h1c2;
						arA23['hc] = 'h15a;
					end
					10: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'h1e3;
						arA23['hc] = 'h15a;
					end
					11: begin
						arIll['hc] = 1'b0;
						arA1['hc] = 'hea;
						arA23['hc] = 'h15b;
					end
					default: begin
						arIll['hc] = 1'b1;
						arA1['hc] = 1'sbx;
						arA23['hc] = 1'sbx;
					end
				endcase
		endcase
		(* full_case, parallel_case *)
		case (row86)
			3'b000:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h1c1;
						arA23['hd] = 1'sbx;
					end
					1: begin
						arIll['hd] = 1'b1;
						arA1['hd] = 1'sbx;
						arA23['hd] = 1'sbx;
					end
					2: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h6;
						arA23['hd] = 'h1c3;
					end
					3: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h21c;
						arA23['hd] = 'h1c3;
					end
					4: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h103;
						arA23['hd] = 'h1c3;
					end
					5: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h1c2;
						arA23['hd] = 'h1c3;
					end
					6: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h1e3;
						arA23['hd] = 'h1c3;
					end
					7: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'ha;
						arA23['hd] = 'h1c3;
					end
					8: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h1e2;
						arA23['hd] = 'h1c3;
					end
					9: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h1c2;
						arA23['hd] = 'h1c3;
					end
					10: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h1e3;
						arA23['hd] = 'h1c3;
					end
					11: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'hea;
						arA23['hd] = 'h1c1;
					end
					default: begin
						arIll['hd] = 1'b1;
						arA1['hd] = 1'sbx;
						arA23['hd] = 1'sbx;
					end
				endcase
			3'b001:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h1c1;
						arA23['hd] = 1'sbx;
					end
					1: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h1c1;
						arA23['hd] = 1'sbx;
					end
					2: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h6;
						arA23['hd] = 'h1c3;
					end
					3: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h21c;
						arA23['hd] = 'h1c3;
					end
					4: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h103;
						arA23['hd] = 'h1c3;
					end
					5: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h1c2;
						arA23['hd] = 'h1c3;
					end
					6: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h1e3;
						arA23['hd] = 'h1c3;
					end
					7: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'ha;
						arA23['hd] = 'h1c3;
					end
					8: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h1e2;
						arA23['hd] = 'h1c3;
					end
					9: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h1c2;
						arA23['hd] = 'h1c3;
					end
					10: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h1e3;
						arA23['hd] = 'h1c3;
					end
					11: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'hea;
						arA23['hd] = 'h1c1;
					end
					default: begin
						arIll['hd] = 1'b1;
						arA1['hd] = 1'sbx;
						arA23['hd] = 1'sbx;
					end
				endcase
			3'b010:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h1c5;
						arA23['hd] = 1'sbx;
					end
					1: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h1c5;
						arA23['hd] = 1'sbx;
					end
					2: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'hb;
						arA23['hd] = 'h1cb;
					end
					3: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'hf;
						arA23['hd] = 'h1cb;
					end
					4: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h179;
						arA23['hd] = 'h1cb;
					end
					5: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h1c6;
						arA23['hd] = 'h1cb;
					end
					6: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h1e7;
						arA23['hd] = 'h1cb;
					end
					7: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'he;
						arA23['hd] = 'h1cb;
					end
					8: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h1e6;
						arA23['hd] = 'h1cb;
					end
					9: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h1c6;
						arA23['hd] = 'h1cb;
					end
					10: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h1e7;
						arA23['hd] = 'h1cb;
					end
					11: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'ha7;
						arA23['hd] = 'h1c5;
					end
					default: begin
						arIll['hd] = 1'b1;
						arA1['hd] = 1'sbx;
						arA23['hd] = 1'sbx;
					end
				endcase
			3'b011:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h1c9;
						arA23['hd] = 1'sbx;
					end
					1: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h1c9;
						arA23['hd] = 1'sbx;
					end
					2: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h6;
						arA23['hd] = 'h1c7;
					end
					3: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h21c;
						arA23['hd] = 'h1c7;
					end
					4: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h103;
						arA23['hd] = 'h1c7;
					end
					5: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h1c2;
						arA23['hd] = 'h1c7;
					end
					6: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h1e3;
						arA23['hd] = 'h1c7;
					end
					7: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'ha;
						arA23['hd] = 'h1c7;
					end
					8: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h1e2;
						arA23['hd] = 'h1c7;
					end
					9: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h1c2;
						arA23['hd] = 'h1c7;
					end
					10: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h1e3;
						arA23['hd] = 'h1c7;
					end
					11: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'hea;
						arA23['hd] = 'h1c9;
					end
					default: begin
						arIll['hd] = 1'b1;
						arA1['hd] = 1'sbx;
						arA23['hd] = 1'sbx;
					end
				endcase
			3'b100:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h1c1;
						arA23['hd] = 1'sbx;
					end
					1: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h10f;
						arA23['hd] = 1'sbx;
					end
					2: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h6;
						arA23['hd] = 'h299;
					end
					3: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h21c;
						arA23['hd] = 'h299;
					end
					4: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h103;
						arA23['hd] = 'h299;
					end
					5: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h1c2;
						arA23['hd] = 'h299;
					end
					6: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h1e3;
						arA23['hd] = 'h299;
					end
					7: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'ha;
						arA23['hd] = 'h299;
					end
					8: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h1e2;
						arA23['hd] = 'h299;
					end
					9: begin
						arIll['hd] = 1'b1;
						arA1['hd] = 1'sbx;
						arA23['hd] = 1'sbx;
					end
					10: begin
						arIll['hd] = 1'b1;
						arA1['hd] = 1'sbx;
						arA23['hd] = 1'sbx;
					end
					11: begin
						arIll['hd] = 1'b1;
						arA1['hd] = 1'sbx;
						arA23['hd] = 1'sbx;
					end
					default: begin
						arIll['hd] = 1'b1;
						arA1['hd] = 1'sbx;
						arA23['hd] = 1'sbx;
					end
				endcase
			3'b101:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h1c1;
						arA23['hd] = 1'sbx;
					end
					1: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h10f;
						arA23['hd] = 1'sbx;
					end
					2: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h6;
						arA23['hd] = 'h299;
					end
					3: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h21c;
						arA23['hd] = 'h299;
					end
					4: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h103;
						arA23['hd] = 'h299;
					end
					5: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h1c2;
						arA23['hd] = 'h299;
					end
					6: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h1e3;
						arA23['hd] = 'h299;
					end
					7: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'ha;
						arA23['hd] = 'h299;
					end
					8: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h1e2;
						arA23['hd] = 'h299;
					end
					9: begin
						arIll['hd] = 1'b1;
						arA1['hd] = 1'sbx;
						arA23['hd] = 1'sbx;
					end
					10: begin
						arIll['hd] = 1'b1;
						arA1['hd] = 1'sbx;
						arA23['hd] = 1'sbx;
					end
					11: begin
						arIll['hd] = 1'b1;
						arA1['hd] = 1'sbx;
						arA23['hd] = 1'sbx;
					end
					default: begin
						arIll['hd] = 1'b1;
						arA1['hd] = 1'sbx;
						arA23['hd] = 1'sbx;
					end
				endcase
			3'b110:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h1c5;
						arA23['hd] = 1'sbx;
					end
					1: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h10b;
						arA23['hd] = 1'sbx;
					end
					2: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'hb;
						arA23['hd] = 'h29d;
					end
					3: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'hf;
						arA23['hd] = 'h29d;
					end
					4: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h179;
						arA23['hd] = 'h29d;
					end
					5: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h1c6;
						arA23['hd] = 'h29d;
					end
					6: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h1e7;
						arA23['hd] = 'h29d;
					end
					7: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'he;
						arA23['hd] = 'h29d;
					end
					8: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h1e6;
						arA23['hd] = 'h29d;
					end
					9: begin
						arIll['hd] = 1'b1;
						arA1['hd] = 1'sbx;
						arA23['hd] = 1'sbx;
					end
					10: begin
						arIll['hd] = 1'b1;
						arA1['hd] = 1'sbx;
						arA23['hd] = 1'sbx;
					end
					11: begin
						arIll['hd] = 1'b1;
						arA1['hd] = 1'sbx;
						arA23['hd] = 1'sbx;
					end
					default: begin
						arIll['hd] = 1'b1;
						arA1['hd] = 1'sbx;
						arA23['hd] = 1'sbx;
					end
				endcase
			3'b111:
				(* full_case, parallel_case *)
				case (col)
					0: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h1c5;
						arA23['hd] = 1'sbx;
					end
					1: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h1c5;
						arA23['hd] = 1'sbx;
					end
					2: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'hb;
						arA23['hd] = 'h1cb;
					end
					3: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'hf;
						arA23['hd] = 'h1cb;
					end
					4: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h179;
						arA23['hd] = 'h1cb;
					end
					5: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h1c6;
						arA23['hd] = 'h1cb;
					end
					6: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h1e7;
						arA23['hd] = 'h1cb;
					end
					7: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'he;
						arA23['hd] = 'h1cb;
					end
					8: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h1e6;
						arA23['hd] = 'h1cb;
					end
					9: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h1c6;
						arA23['hd] = 'h1cb;
					end
					10: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'h1e7;
						arA23['hd] = 'h1cb;
					end
					11: begin
						arIll['hd] = 1'b0;
						arA1['hd] = 'ha7;
						arA23['hd] = 'h1c5;
					end
					default: begin
						arIll['hd] = 1'b1;
						arA1['hd] = 1'sbx;
						arA23['hd] = 1'sbx;
					end
				endcase
		endcase
	end
	initial _sv2v_0 = 0;
endmodule
